magic
tech sky130A
magscale 1 2
timestamp 1744462317
<< locali >>
rect 2048 -7782 2240 -7264
rect 2048 -7962 2054 -7782
rect 2234 -7962 2240 -7782
rect 2048 -7968 2240 -7962
<< viali >>
rect 3360 -7424 3552 -7232
rect 2054 -7962 2234 -7782
<< metal1 >>
rect 2048 -7782 2240 -7770
rect 2048 -7962 2054 -7782
rect 2234 -7962 2240 -7782
rect 2048 -8704 2240 -7962
rect 2304 -8256 2496 -4096
rect 3348 -7232 3564 -7226
rect 3348 -7424 3360 -7232
rect 3552 -7424 3564 -7232
rect 3348 -7430 3564 -7424
rect 3360 -7456 3552 -7430
rect 3360 -7654 3552 -7648
rect 1920 -9184 1984 -8800
rect 2304 -9248 2496 -8728
rect 2304 -9440 2528 -9248
rect 2720 -9440 2726 -9248
<< via1 >>
rect 3360 -7648 3552 -7456
rect 2528 -9440 2720 -9248
<< metal2 >>
rect 3354 -7648 3360 -7456
rect 3552 -7648 3558 -7456
rect 3360 -7712 3552 -7648
rect 3360 -7913 3552 -7904
rect 2528 -9248 2720 -9242
rect 2784 -9248 2976 -9239
rect 2720 -9440 2784 -9248
rect 2528 -9446 2720 -9440
rect 2784 -9449 2976 -9440
<< via2 >>
rect 3360 -7904 3552 -7712
rect 2784 -9440 2976 -9248
<< metal3 >>
rect 3355 -7712 3557 -7707
rect 3355 -7904 3360 -7712
rect 3552 -7904 3557 -7712
rect 3355 -7909 3557 -7904
rect 3360 -8032 3552 -7909
rect 3360 -8230 3552 -8224
rect 2779 -9248 2981 -9243
rect 2779 -9440 2784 -9248
rect 2976 -9440 2981 -9248
rect 2779 -9445 2981 -9440
rect 2784 -9792 2977 -9445
rect -3200 -9920 8576 -9792
rect 2784 -9952 2977 -9920
rect 8024 -12790 8124 -10004
rect -3176 -12890 8524 -12790
rect 8024 -15890 8124 -12890
rect -3176 -15990 8524 -15890
rect 8024 -18890 8124 -15990
rect -3176 -18990 8524 -18890
rect 8024 -21990 8124 -18990
rect -3176 -22090 8524 -21990
rect 8024 -24490 8124 -22090
<< via3 >>
rect 3360 -8224 3552 -8032
<< metal4 >>
rect 3359 -8032 3553 -8031
rect 3359 -8224 3360 -8032
rect 3552 -8224 3553 -8032
rect 3359 -8225 3553 -8224
rect 3360 -9792 3552 -8225
rect -3200 -9920 3012 -9792
rect 3220 -9920 8576 -9792
rect 3360 -10016 3552 -9920
rect 8024 -12790 8124 -9940
rect -3176 -12890 8524 -12790
rect 8024 -15890 8124 -12890
rect -3176 -15990 8524 -15890
rect 8024 -18890 8124 -15990
rect -3176 -18990 8524 -18890
rect 8024 -21990 8124 -18990
rect -3176 -22090 8524 -21990
rect 8024 -24490 8124 -22090
use JNWTR_CAPX4  x1_0 ../JNW_TR_SKY130A
timestamp 1744451459
transform -1 0 2956 0 -1 -9786
box 480 0 3120 2640
use JNWTR_CAPX4  x1_1
timestamp 1744451459
transform -1 0 2956 0 -1 -12826
box 480 0 3120 2640
use JNWTR_CAPX4  x1_2
timestamp 1744451459
transform -1 0 2956 0 -1 -15866
box 480 0 3120 2640
use JNWTR_CAPX4  x1_3
timestamp 1744451459
transform -1 0 2956 0 -1 -18906
box 480 0 3120 2640
use JNWTR_CAPX4  x1_4
timestamp 1744451459
transform -1 0 2956 0 -1 -21946
box 480 0 3120 2640
use JNWTR_CAPX4  x1_5
timestamp 1744451459
transform -1 0 9056 0 -1 -9786
box 480 0 3120 2640
use JNWTR_CAPX4  x1_6
timestamp 1744451459
transform -1 0 9056 0 -1 -12826
box 480 0 3120 2640
use JNWTR_CAPX4  x1_7
timestamp 1744451459
transform 1 0 5456 0 -1 -15866
box 480 0 3120 2640
use JNWTR_CAPX4  x1_8
timestamp 1744451459
transform -1 0 9056 0 -1 -18906
box 480 0 3120 2640
use JNWTR_CAPX4  x1_9
timestamp 1744451459
transform -1 0 9056 0 -1 -21946
box 480 0 3120 2640
use JNWTR_CAPX4  x1_10
timestamp 1744451459
transform -1 0 -76 0 -1 -9790
box 480 0 3120 2640
use JNWTR_CAPX4  x1_11
timestamp 1744451459
transform -1 0 -76 0 -1 -12830
box 480 0 3120 2640
use JNWTR_CAPX4  x1_12
timestamp 1744451459
transform -1 0 -76 0 -1 -15870
box 480 0 3120 2640
use JNWTR_CAPX4  x1_13
timestamp 1744451459
transform -1 0 -76 0 -1 -18910
box 480 0 3120 2640
use JNWTR_CAPX4  x1_14
timestamp 1744451459
transform -1 0 -76 0 -1 -21950
box 480 0 3120 2640
use JNWTR_CAPX4  x1_15
timestamp 1744451459
transform -1 0 6024 0 -1 -9790
box 480 0 3120 2640
use JNWTR_CAPX4  x1_16
timestamp 1744451459
transform -1 0 6024 0 -1 -12830
box 480 0 3120 2640
use JNWTR_CAPX4  x1_17
timestamp 1744451459
transform -1 0 6024 0 -1 -15870
box 480 0 3120 2640
use JNWTR_CAPX4  x1_18
timestamp 1744451459
transform -1 0 6024 0 -1 -18910
box 480 0 3120 2640
use JNWTR_CAPX4  x1_19
timestamp 1744451459
transform -1 0 6024 0 -1 -21950
box 480 0 3120 2640
use JNWATR_NCH_2C5F0  x4 ../JNW_ATR_SKY130A
timestamp 1744458479
transform 1 0 1760 0 -1 -8160
box -184 -128 1208 928
use JNW_VIS_OTA  x7 ../JNW_GR02_SKY130A
timestamp 1744462317
transform 1 0 4768 0 1 -4648
box -9120 -3400 4936 2656
<< labels >>
flabel metal1 2304 -9408 2496 -9216 0 FreeSans 400 0 0 0 I_TEMP
flabel metal1 1920 -9184 1984 -9120 0 FreeSans 400 0 0 0 DISCHARGE
<< properties >>
string FIXED_BBOX 0 0 6008 7240
<< end >>
