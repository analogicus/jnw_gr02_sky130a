magic
tech sky130A
magscale 1 2
timestamp 1744464884
<< metal1 >>
rect 18976 6501 19488 6693
rect -14100 4892 -1456 5084
rect 988 3636 2854 3700
rect 3732 3232 3924 5744
rect 19296 4960 19488 6501
rect 14560 4768 19488 4960
rect 3732 3040 12000 3232
<< metal3 >>
rect 15848 4480 18520 4608
rect 15308 3136 15484 3960
rect 15848 3704 16024 4480
rect 17804 3136 17980 4024
rect 18344 3704 18520 4480
rect 15308 3008 17984 3136
use JNW_VIS_ITIME  x1 ../JNW_GR02_SKY130A
timestamp 1744463149
transform 1 0 9521 0 1 12525
box -4352 -24590 9981 -1992
use JNW_VIS_TI  x2 ../JNW_GR02_SKY130A
timestamp 1744464884
transform 1 0 -5504 0 1 13448
box -9344 -19400 9900 -2398
use JNWTR_DFTSPCX1_CV  x3 ../JNW_TR_SKY130A
timestamp 1744464884
transform 1 0 14678 0 1 3320
box -150 -120 2130 1080
use JNWTR_DFTSPCX1_CV  x4
timestamp 1744464884
transform 1 0 17174 0 1 3320
box -150 -120 2130 1080
use dig  x5 ../JNW_GR02_SKY130A
timestamp 1744463149
transform 1 0 -10247 0 1 -20067
box 0 824 9395 10464
<< properties >>
string FIXED_BBOX 0 0 22267 11539
<< end >>
