.subckt dig VGND VPWR clk counter_out[0] counter_out[1] counter_out[2] counter_out[3]
+ counter_out[4] counter_out[5] counter_out[6] counter_out[7] trigger
XTAP_TAPCELL_ROW_26_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_49_ net25 _25_ _16_ VGND VGND VPWR VPWR _28_ sky130_fd_sc_hd__o21ai_1
X_66_ clknet_1_1__leaf_clk _04_ VGND VGND VPWR VPWR counter\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_17_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput7 net7 VGND VGND VPWR VPWR counter_out[5] sky130_fd_sc_hd__buf_2
XFILLER_3_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_65_ clknet_1_0__leaf_clk _03_ VGND VGND VPWR VPWR counter\[3\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Left_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_48_ counter\[4\] counter\[5\] counter\[6\] _21_ VGND VGND VPWR VPWR _27_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_12_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput8 net8 VGND VGND VPWR VPWR counter_out[6] sky130_fd_sc_hd__buf_2
XFILLER_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_47_ _25_ _26_ VGND VGND VPWR VPWR _05_ sky130_fd_sc_hd__nor2_1
X_64_ clknet_1_0__leaf_clk _02_ VGND VGND VPWR VPWR counter\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold10 net6 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput9 net9 VGND VGND VPWR VPWR counter_out[7] sky130_fd_sc_hd__buf_2
XFILLER_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_63_ clknet_1_0__leaf_clk _01_ VGND VGND VPWR VPWR counter\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_46_ _16_ _24_ VGND VGND VPWR VPWR _26_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold11 _12_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_62_ clknet_1_0__leaf_clk _00_ VGND VGND VPWR VPWR counter\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_34_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold12 net7 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlygate4sd3_1
X_45_ counter\[4\] counter\[5\] _21_ VGND VGND VPWR VPWR _25_ sky130_fd_sc_hd__and3_1
XFILLER_18_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload0 clknet_1_0__leaf_clk VGND VGND VPWR VPWR clkload0/X sky130_fd_sc_hd__clkbuf_4
XFILLER_31_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_61_ counter\[7\] net16 _30_ VGND VGND VPWR VPWR _15_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_19_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_44_ counter\[4\] _21_ counter\[5\] VGND VGND VPWR VPWR _24_ sky130_fd_sc_hd__a21o_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold13 _13_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_60_ counter\[6\] net14 _30_ VGND VGND VPWR VPWR _14_ sky130_fd_sc_hd__mux2_1
XFILLER_23_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_20_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_43_ net26 _21_ _23_ VGND VGND VPWR VPWR _04_ sky130_fd_sc_hd__a21oi_1
Xhold14 net2 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_35_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_42_ counter\[4\] _21_ _16_ VGND VGND VPWR VPWR _23_ sky130_fd_sc_hd__o21ai_1
Xhold15 counter\[7\] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_41_ _16_ _20_ _22_ VGND VGND VPWR VPWR _03_ sky130_fd_sc_hd__and3_1
XFILLER_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold16 counter\[6\] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_40_ _21_ VGND VGND VPWR VPWR _22_ sky130_fd_sc_hd__inv_2
Xhold17 counter\[4\] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_27_Left_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_11_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput1 trigger VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_10_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_78_ clknet_1_1__leaf_clk net1 VGND VGND VPWR VPWR trigger_prev sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_77_ clknet_1_1__leaf_clk net17 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dfxtp_1
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_76_ clknet_1_1__leaf_clk net15 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dfxtp_1
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_59_ counter\[5\] net21 _30_ VGND VGND VPWR VPWR _13_ sky130_fd_sc_hd__mux2_1
XFILLER_7_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_23_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_75_ clknet_1_1__leaf_clk net22 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dfxtp_1
X_58_ counter\[4\] net19 _30_ VGND VGND VPWR VPWR _12_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Left_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_74_ clknet_1_1__leaf_clk net20 VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dfxtp_1
XFILLER_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_57_ counter\[3\] net12 _30_ VGND VGND VPWR VPWR _11_ sky130_fd_sc_hd__mux2_1
XFILLER_27_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_73_ clknet_1_0__leaf_clk net13 VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dfxtp_1
X_56_ counter\[2\] net10 _30_ VGND VGND VPWR VPWR _10_ sky130_fd_sc_hd__mux2_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_39_ counter\[0\] counter\[1\] counter\[2\] counter\[3\] VGND VGND VPWR VPWR _21_
+ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_4_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_72_ clknet_1_0__leaf_clk net11 VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dfxtp_1
XFILLER_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_55_ counter\[1\] net18 _30_ VGND VGND VPWR VPWR _09_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_38_ counter\[0\] counter\[1\] counter\[2\] counter\[3\] VGND VGND VPWR VPWR _20_
+ sky130_fd_sc_hd__a31o_1
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1 net4 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_2_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_71_ clknet_1_0__leaf_clk _09_ VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dfxtp_1
X_54_ counter\[0\] net23 _30_ VGND VGND VPWR VPWR _08_ sky130_fd_sc_hd__mux2_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_37_ _16_ _18_ _19_ VGND VGND VPWR VPWR _02_ sky130_fd_sc_hd__and3_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_31_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2 _10_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_34_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_70_ clknet_1_0__leaf_clk _08_ VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dfxtp_1
XFILLER_35_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_53_ trigger_prev net1 VGND VGND VPWR VPWR _30_ sky130_fd_sc_hd__nand2b_4
XFILLER_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36_ counter\[0\] counter\[1\] counter\[2\] VGND VGND VPWR VPWR _19_ sky130_fd_sc_hd__nand3_1
XFILLER_8_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3 net5 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_52_ net24 _27_ _29_ VGND VGND VPWR VPWR _07_ sky130_fd_sc_hd__o21a_1
X_35_ counter\[0\] counter\[1\] counter\[2\] VGND VGND VPWR VPWR _18_ sky130_fd_sc_hd__a21o_1
Xhold4 _11_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_51_ net24 _27_ _16_ VGND VGND VPWR VPWR _29_ sky130_fd_sc_hd__a21boi_1
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34_ counter\[0\] counter\[1\] _17_ VGND VGND VPWR VPWR _01_ sky130_fd_sc_hd__o21a_1
Xhold5 net8 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_50_ _27_ _28_ VGND VGND VPWR VPWR _06_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_22_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33_ counter\[0\] counter\[1\] _16_ VGND VGND VPWR VPWR _17_ sky130_fd_sc_hd__a21boi_1
Xhold6 _14_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_25_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32_ counter\[0\] _16_ VGND VGND VPWR VPWR _00_ sky130_fd_sc_hd__and2b_1
Xhold7 net9 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31_ net1 trigger_prev VGND VGND VPWR VPWR _16_ sky130_fd_sc_hd__nand2b_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold8 _15_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_8_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_29_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold9 net3 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_1_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_30_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_4_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput2 net2 VGND VGND VPWR VPWR counter_out[0] sky130_fd_sc_hd__buf_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput3 net3 VGND VGND VPWR VPWR counter_out[1] sky130_fd_sc_hd__buf_2
X_69_ clknet_1_1__leaf_clk _07_ VGND VGND VPWR VPWR counter\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_8_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput4 net4 VGND VGND VPWR VPWR counter_out[2] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_68_ clknet_1_1__leaf_clk _06_ VGND VGND VPWR VPWR counter\[6\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_24_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput5 net5 VGND VGND VPWR VPWR counter_out[3] sky130_fd_sc_hd__buf_2
XFILLER_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_67_ clknet_1_1__leaf_clk _05_ VGND VGND VPWR VPWR counter\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput6 net6 VGND VGND VPWR VPWR counter_out[4] sky130_fd_sc_hd__buf_2
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
.ends

