** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_GR02_SKY130A/JNW_VIS_TI.sch
.subckt JNW_VIS_TI I_TEMP VDD VREF LPO LPI PWR_UP VSS
*.ipin VSS
*.opin VREF
*.ipin PWR_UP
*.opin LPI
*.opin LPO
*.ipin VDD
*.opin I_TEMP
XQ1 VSS VSS VIN sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1 mult=1
XQ2 VSS VSS VD2 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=8 mult=8
x7 VDD VIN VIP VSS LPO JNW_VIS_OTA
x11 LPI PWR_UP VSS VSS JNWATR_NCH_12C5F0
x1<0> LPI VSS JNWTR_CAPX4
x1<1> LPI VSS JNWTR_CAPX4
x1<2> LPI VSS JNWTR_CAPX4
x1<3> LPI VSS JNWTR_CAPX4
x9 V_MEAS1 LPI VSS VSS JNWATR_NCH_12C5F0
x2<0> V_MEAS2 V_MEAS1 VDD VDD JNWATR_PCH_4C5F0
x2<1> V_MEAS2 V_MEAS1 VDD VDD JNWATR_PCH_4C5F0
x2<2> V_MEAS2 V_MEAS1 VDD VDD JNWATR_PCH_4C5F0
x3<0> V_MEAS1 V_MEAS3 V_MEAS2 V_MEAS2 JNWATR_PCH_4C5F0
x3<1> V_MEAS1 V_MEAS3 V_MEAS2 V_MEAS2 JNWATR_PCH_4C5F0
x3<2> V_MEAS1 V_MEAS3 V_MEAS2 V_MEAS2 JNWATR_PCH_4C5F0
x4<0> V_MEAS4 V_MEAS1 VDD VDD JNWATR_PCH_4C5F0
x4<1> V_MEAS4 V_MEAS1 VDD VDD JNWATR_PCH_4C5F0
x4<2> V_MEAS4 V_MEAS1 VDD VDD JNWATR_PCH_4C5F0
x5<0> VREF V_MEAS3 V_MEAS4 V_MEAS4 JNWATR_PCH_4C5F0
x5<1> VREF V_MEAS3 V_MEAS4 V_MEAS4 JNWATR_PCH_4C5F0
x5<2> VREF V_MEAS3 V_MEAS4 V_MEAS4 JNWATR_PCH_4C5F0
x15 V_MEAS3 V_MEAS3 VDD VDD JNWATR_PCH_2C5F0
x7<0> V_MEAS5 V_MEAS1 VDD VDD JNWATR_PCH_4C5F0
x7<1> V_MEAS5 V_MEAS1 VDD VDD JNWATR_PCH_4C5F0
x7<2> V_MEAS5 V_MEAS1 VDD VDD JNWATR_PCH_4C5F0
xa1<0> VIN V_MEAS3 V_MEAS5 V_MEAS5 JNWATR_PCH_4C5F0
xa1<1> VIN V_MEAS3 V_MEAS5 V_MEAS5 JNWATR_PCH_4C5F0
xa1<2> VIN V_MEAS3 V_MEAS5 V_MEAS5 JNWATR_PCH_4C5F0
x14 VIP VREF VSS JNWTR_RPPO4
x13<0> VD2 VIP VSS JNWTR_RPPO2
x13<1> VD2 VIP VSS JNWTR_RPPO2
x13<2> VD2 VIP VSS JNWTR_RPPO2
x13<3> VD2 VIP VSS JNWTR_RPPO2
x3 VSS V_MEAS3 VSS JNWTR_RPPO2
x2 V_MEAS6 V_MEAS1 VDD VDD JNWATR_PCH_2C5F0
x16<0> I_TEMP V_MEAS3 V_MEAS6 V_MEAS6 JNWATR_PCH_4C5F0
x16<1> I_TEMP V_MEAS3 V_MEAS6 V_MEAS6 JNWATR_PCH_4C5F0
x16<2> I_TEMP V_MEAS3 V_MEAS6 V_MEAS6 JNWATR_PCH_4C5F0
.ends

* expanding   symbol:  JNW_GR02_SKY130A/JNW_VIS_OTA.sym # of pins=5
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_GR02_SKY130A/JNW_VIS_OTA.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_GR02_SKY130A/JNW_VIS_OTA.sch
.subckt JNW_VIS_OTA VDD VIN VIP VSS VOUT
*.ipin VDD
*.ipin VIP
*.ipin VIN
*.ipin VSS
*.opin VOUT
xd01<0> V2 VIP VOP VDD JNWATR_PCH_12C1F2
xd01<1> V2 VIP VOP VDD JNWATR_PCH_12C1F2
xd01<2> V2 VIP VOP VDD JNWATR_PCH_12C1F2
xd01<3> V2 VIP VOP VDD JNWATR_PCH_12C1F2
xd02<0> V1 VIN VOP VDD JNWATR_PCH_12C1F2
xd02<1> V1 VIN VOP VDD JNWATR_PCH_12C1F2
xd02<2> V1 VIN VOP VDD JNWATR_PCH_12C1F2
xd02<3> V1 VIN VOP VDD JNWATR_PCH_12C1F2
xc04 VOUT V1 VSS VSS JNWATR_NCH_12C5F0
xc02 V2 V2 VSS VSS JNWATR_NCH_12C5F0
xc01 net1 V2 VSS VSS JNWATR_NCH_12C5F0
xc03 V1 V1 VSS VSS JNWATR_NCH_12C5F0
xb02<0> VOUT net1 VDD VDD JNWATR_PCH_12C5F0
xb02<1> VOUT net1 VDD VDD JNWATR_PCH_12C5F0
xb02<2> VOUT net1 VDD VDD JNWATR_PCH_12C5F0
xb02<3> VOUT net1 VDD VDD JNWATR_PCH_12C5F0
xb01<0> net1 net1 VDD VDD JNWATR_PCH_12C5F0
xb01<1> net1 net1 VDD VDD JNWATR_PCH_12C5F0
xb01<2> net1 net1 VDD VDD JNWATR_PCH_12C5F0
xb01<3> net1 net1 VDD VDD JNWATR_PCH_12C5F0
x6 net3 net2 VSS JNWTR_RPPO2
x8<0> VSS net3 VSS JNWTR_RPPO2
x8<1> VSS net3 VSS JNWTR_RPPO2
xa01 net2 net2 VDD VDD JNWATR_PCH_12C5F0
xa02 VOP net2 VDD VDD JNWATR_PCH_12C5F0
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_12C5F0.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_12C5F0.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_12C5F0.sch
.subckt JNWATR_NCH_12C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.94 W=8.32 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_CAPX4.sym # of pins=2
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX4.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX4.sch
.subckt JNWTR_CAPX4 A B
*.iopin A
*.iopin B
XXA1 A B JNWTR_CAPX1
XXA2 A B JNWTR_CAPX1
XXB1 A B JNWTR_CAPX1
XXB2 A B JNWTR_CAPX1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sch
.subckt JNWATR_PCH_4C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.94 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_2C5F0.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_2C5F0.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_2C5F0.sch
.subckt JNWATR_PCH_2C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.94 W=1.92 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RPPO4.sym # of pins=3
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO4.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO4.sch
.subckt JNWTR_RPPO4 N P B
*.iopin P
*.iopin N
*.iopin B
XXA1 N P B JNWTR_RES4
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RPPO2.sym # of pins=3
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO2.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO2.sch
.subckt JNWTR_RPPO2 N P B
*.iopin P
*.iopin N
*.iopin B
XXA1 N P B JNWTR_RES2
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_12C1F2.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_12C1F2.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_12C1F2.sch
.subckt JNWATR_PCH_12C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.22 W=8.32 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_12C5F0.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_12C5F0.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_12C5F0.sch
.subckt JNWATR_PCH_12C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.94 W=8.32 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_CAPX1.sym # of pins=2
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sch
.subckt JNWTR_CAPX1 A B
*.iopin A
*.iopin B
XC1 B A sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RES4.sym # of pins=3
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RES4.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RES4.sch
.subckt JNWTR_RES4 N P B
*.iopin N
*.iopin P
*.iopin B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_1 INT_1 INT_0 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_2 INT_2 INT_1 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_3 P INT_2 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RES2.sym # of pins=3
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RES2.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RES2.sch
.subckt JNWTR_RES2 N P B
*.iopin N
*.iopin P
*.iopin B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_1 P INT_0 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
.ends

.end
