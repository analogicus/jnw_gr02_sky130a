magic
tech sky130A
magscale 1 2
timestamp 1744552703
<< viali >>
rect 4997 21641 5031 21675
rect 4813 21505 4847 21539
rect 4997 20961 5031 20995
rect 4445 20757 4479 20791
rect 5089 20553 5123 20587
rect 2237 20417 2271 20451
rect 2504 20417 2538 20451
rect 3709 20417 3743 20451
rect 3976 20417 4010 20451
rect 3617 20213 3651 20247
rect 2421 20009 2455 20043
rect 3617 19873 3651 19907
rect 4721 19873 4755 19907
rect 2605 19805 2639 19839
rect 2789 19805 2823 19839
rect 2881 19805 2915 19839
rect 2973 19805 3007 19839
rect 4445 19805 4479 19839
rect 4537 19737 4571 19771
rect 4077 19669 4111 19703
rect 2881 19465 2915 19499
rect 2973 19465 3007 19499
rect 4077 19465 4111 19499
rect 4997 19465 5031 19499
rect 2789 19329 2823 19363
rect 4813 19329 4847 19363
rect 3249 19261 3283 19295
rect 4629 19261 4663 19295
rect 2329 18921 2363 18955
rect 1961 18717 1995 18751
rect 2421 18717 2455 18751
rect 4721 18717 4755 18751
rect 4077 18581 4111 18615
rect 2789 18377 2823 18411
rect 5089 18377 5123 18411
rect 3976 18309 4010 18343
rect 1409 18241 1443 18275
rect 1676 18241 1710 18275
rect 3709 18241 3743 18275
rect 3065 18173 3099 18207
rect 3617 18037 3651 18071
rect 4169 17833 4203 17867
rect 1593 17765 1627 17799
rect 2697 17765 2731 17799
rect 4629 17697 4663 17731
rect 4813 17697 4847 17731
rect 1409 17629 1443 17663
rect 2237 17629 2271 17663
rect 3157 17629 3191 17663
rect 4537 17493 4571 17527
rect 3065 17153 3099 17187
rect 3332 17153 3366 17187
rect 4445 16949 4479 16983
rect 2973 16745 3007 16779
rect 3341 16745 3375 16779
rect 2881 16677 2915 16711
rect 2789 16609 2823 16643
rect 4353 16609 4387 16643
rect 3065 16541 3099 16575
rect 3157 16541 3191 16575
rect 3341 16541 3375 16575
rect 4813 16541 4847 16575
rect 3801 16473 3835 16507
rect 4997 16405 5031 16439
rect 2053 16065 2087 16099
rect 2237 16065 2271 16099
rect 2053 15861 2087 15895
rect 2973 15657 3007 15691
rect 1409 15453 1443 15487
rect 4629 15453 4663 15487
rect 1676 15385 1710 15419
rect 3157 15385 3191 15419
rect 3249 15385 3283 15419
rect 3525 15385 3559 15419
rect 2789 15317 2823 15351
rect 3341 15317 3375 15351
rect 4077 15317 4111 15351
rect 1961 15113 1995 15147
rect 2513 15113 2547 15147
rect 2145 15045 2179 15079
rect 1869 14977 1903 15011
rect 2053 14977 2087 15011
rect 2329 14977 2363 15011
rect 2605 14977 2639 15011
rect 2697 14977 2731 15011
rect 3985 14773 4019 14807
rect 2513 14569 2547 14603
rect 2697 14569 2731 14603
rect 4077 14569 4111 14603
rect 4721 14433 4755 14467
rect 3065 14365 3099 14399
rect 4445 14365 4479 14399
rect 2665 14297 2699 14331
rect 2881 14297 2915 14331
rect 3617 14297 3651 14331
rect 4537 14297 4571 14331
rect 5089 14025 5123 14059
rect 3976 13957 4010 13991
rect 3709 13821 3743 13855
rect 3801 13413 3835 13447
rect 4905 13413 4939 13447
rect 3157 13345 3191 13379
rect 4445 13345 4479 13379
rect 4169 13277 4203 13311
rect 5089 13277 5123 13311
rect 2605 13141 2639 13175
rect 4261 13141 4295 13175
rect 2237 12937 2271 12971
rect 4445 12937 4479 12971
rect 2421 12869 2455 12903
rect 2145 12801 2179 12835
rect 2605 12801 2639 12835
rect 4997 12733 5031 12767
rect 2421 12597 2455 12631
rect 3893 12597 3927 12631
rect 3065 12393 3099 12427
rect 2973 12257 3007 12291
rect 4537 12257 4571 12291
rect 1501 12189 1535 12223
rect 3157 12189 3191 12223
rect 3249 12189 3283 12223
rect 1768 12121 1802 12155
rect 2881 12053 2915 12087
rect 3893 12053 3927 12087
rect 4997 11849 5031 11883
rect 2205 11781 2239 11815
rect 2421 11781 2455 11815
rect 3884 11781 3918 11815
rect 3617 11713 3651 11747
rect 2053 11509 2087 11543
rect 2237 11509 2271 11543
rect 1593 11305 1627 11339
rect 4169 11237 4203 11271
rect 1685 11101 1719 11135
rect 1777 11101 1811 11135
rect 2044 11101 2078 11135
rect 4353 11101 4387 11135
rect 5089 11101 5123 11135
rect 3157 10965 3191 10999
rect 4445 10965 4479 10999
rect 2329 10761 2363 10795
rect 5089 10761 5123 10795
rect 3617 10693 3651 10727
rect 3954 10693 3988 10727
rect 3709 10625 3743 10659
rect 2513 10557 2547 10591
rect 2605 10557 2639 10591
rect 2697 10557 2731 10591
rect 2789 10557 2823 10591
rect 3065 10557 3099 10591
rect 4077 10217 4111 10251
rect 3065 10081 3099 10115
rect 4721 10081 4755 10115
rect 3249 10013 3283 10047
rect 4445 10013 4479 10047
rect 2513 9945 2547 9979
rect 3617 9945 3651 9979
rect 4537 9945 4571 9979
rect 3341 9877 3375 9911
rect 3433 9877 3467 9911
rect 3985 9673 4019 9707
rect 2697 9605 2731 9639
rect 2145 9537 2179 9571
rect 2237 9537 2271 9571
rect 2421 9537 2455 9571
rect 2605 9333 2639 9367
rect 3065 9129 3099 9163
rect 2789 9061 2823 9095
rect 1409 8925 1443 8959
rect 3341 8925 3375 8959
rect 5089 8925 5123 8959
rect 1676 8857 1710 8891
rect 3249 8857 3283 8891
rect 3433 8857 3467 8891
rect 3617 8857 3651 8891
rect 2881 8789 2915 8823
rect 3049 8789 3083 8823
rect 3341 8789 3375 8823
rect 4445 8789 4479 8823
rect 5089 8585 5123 8619
rect 3617 8517 3651 8551
rect 3954 8517 3988 8551
rect 3709 8449 3743 8483
rect 3065 8381 3099 8415
rect 3985 8041 4019 8075
rect 4537 7905 4571 7939
rect 4353 7837 4387 7871
rect 4445 7837 4479 7871
rect 4813 7837 4847 7871
rect 4997 7701 5031 7735
rect 3065 7293 3099 7327
rect 3341 7225 3375 7259
rect 3525 7157 3559 7191
rect 1409 6817 1443 6851
rect 3341 6817 3375 6851
rect 2881 6749 2915 6783
rect 1676 6681 1710 6715
rect 2973 6681 3007 6715
rect 2789 6613 2823 6647
rect 3065 6613 3099 6647
rect 2053 6409 2087 6443
rect 3678 6341 3712 6375
rect 2237 6273 2271 6307
rect 3433 6273 3467 6307
rect 2513 6205 2547 6239
rect 2421 6137 2455 6171
rect 4813 6069 4847 6103
rect 3617 5661 3651 5695
rect 5089 5661 5123 5695
rect 2973 5525 3007 5559
rect 4445 5525 4479 5559
rect 3249 5321 3283 5355
rect 3157 5185 3191 5219
rect 3709 5185 3743 5219
rect 3976 5185 4010 5219
rect 3433 5117 3467 5151
rect 2789 4981 2823 5015
rect 5089 4981 5123 5015
rect 4261 4777 4295 4811
rect 4721 4641 4755 4675
rect 4813 4641 4847 4675
rect 2237 4573 2271 4607
rect 4629 4573 4663 4607
rect 2504 4505 2538 4539
rect 3617 4437 3651 4471
rect 4813 4097 4847 4131
rect 4997 3961 5031 3995
rect 5089 2397 5123 2431
rect 4905 2261 4939 2295
<< metal1 >>
rect 1104 21786 5428 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 5428 21786
rect 1104 21712 5428 21734
rect 4985 21675 5043 21681
rect 4985 21641 4997 21675
rect 5031 21672 5043 21675
rect 5258 21672 5264 21684
rect 5031 21644 5264 21672
rect 5031 21641 5043 21644
rect 4985 21635 5043 21641
rect 5258 21632 5264 21644
rect 5316 21632 5322 21684
rect 4798 21496 4804 21548
rect 4856 21496 4862 21548
rect 1104 21242 5428 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 5428 21242
rect 1104 21168 5428 21190
rect 4798 20952 4804 21004
rect 4856 20992 4862 21004
rect 4985 20995 5043 21001
rect 4985 20992 4997 20995
rect 4856 20964 4997 20992
rect 4856 20952 4862 20964
rect 4985 20961 4997 20964
rect 5031 20961 5043 20995
rect 4985 20955 5043 20961
rect 4433 20791 4491 20797
rect 4433 20757 4445 20791
rect 4479 20788 4491 20791
rect 4614 20788 4620 20800
rect 4479 20760 4620 20788
rect 4479 20757 4491 20760
rect 4433 20751 4491 20757
rect 4614 20748 4620 20760
rect 4672 20748 4678 20800
rect 1104 20698 5428 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 5428 20698
rect 1104 20624 5428 20646
rect 4798 20544 4804 20596
rect 4856 20584 4862 20596
rect 5077 20587 5135 20593
rect 5077 20584 5089 20587
rect 4856 20556 5089 20584
rect 4856 20544 4862 20556
rect 5077 20553 5089 20556
rect 5123 20553 5135 20587
rect 5077 20547 5135 20553
rect 2240 20488 3740 20516
rect 2240 20457 2268 20488
rect 3712 20460 3740 20488
rect 2498 20457 2504 20460
rect 2225 20451 2283 20457
rect 2225 20417 2237 20451
rect 2271 20417 2283 20451
rect 2225 20411 2283 20417
rect 2492 20411 2504 20457
rect 2498 20408 2504 20411
rect 2556 20408 2562 20460
rect 3694 20408 3700 20460
rect 3752 20408 3758 20460
rect 3970 20457 3976 20460
rect 3964 20411 3976 20457
rect 3970 20408 3976 20411
rect 4028 20408 4034 20460
rect 3602 20204 3608 20256
rect 3660 20204 3666 20256
rect 1104 20154 5428 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 5428 20154
rect 1104 20080 5428 20102
rect 2409 20043 2467 20049
rect 2409 20009 2421 20043
rect 2455 20040 2467 20043
rect 2498 20040 2504 20052
rect 2455 20012 2504 20040
rect 2455 20009 2467 20012
rect 2409 20003 2467 20009
rect 2498 20000 2504 20012
rect 2556 20000 2562 20052
rect 3602 19864 3608 19916
rect 3660 19904 3666 19916
rect 4709 19907 4767 19913
rect 3660 19876 4476 19904
rect 3660 19864 3666 19876
rect 2593 19839 2651 19845
rect 2593 19805 2605 19839
rect 2639 19805 2651 19839
rect 2593 19799 2651 19805
rect 2608 19700 2636 19799
rect 2774 19796 2780 19848
rect 2832 19796 2838 19848
rect 2866 19796 2872 19848
rect 2924 19836 2930 19848
rect 4448 19845 4476 19876
rect 4709 19873 4721 19907
rect 4755 19904 4767 19907
rect 5258 19904 5264 19916
rect 4755 19876 5264 19904
rect 4755 19873 4767 19876
rect 4709 19867 4767 19873
rect 5258 19864 5264 19876
rect 5316 19864 5322 19916
rect 2961 19839 3019 19845
rect 2961 19836 2973 19839
rect 2924 19808 2973 19836
rect 2924 19796 2930 19808
rect 2961 19805 2973 19808
rect 3007 19805 3019 19839
rect 2961 19799 3019 19805
rect 4433 19839 4491 19845
rect 4433 19805 4445 19839
rect 4479 19805 4491 19839
rect 4433 19799 4491 19805
rect 4525 19771 4583 19777
rect 4525 19737 4537 19771
rect 4571 19768 4583 19771
rect 4614 19768 4620 19780
rect 4571 19740 4620 19768
rect 4571 19737 4583 19740
rect 4525 19731 4583 19737
rect 4614 19728 4620 19740
rect 4672 19728 4678 19780
rect 2958 19700 2964 19712
rect 2608 19672 2964 19700
rect 2958 19660 2964 19672
rect 3016 19660 3022 19712
rect 4065 19703 4123 19709
rect 4065 19669 4077 19703
rect 4111 19700 4123 19703
rect 4338 19700 4344 19712
rect 4111 19672 4344 19700
rect 4111 19669 4123 19672
rect 4065 19663 4123 19669
rect 4338 19660 4344 19672
rect 4396 19660 4402 19712
rect 1104 19610 5428 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 5428 19610
rect 1104 19536 5428 19558
rect 2866 19456 2872 19508
rect 2924 19456 2930 19508
rect 2958 19456 2964 19508
rect 3016 19456 3022 19508
rect 3970 19456 3976 19508
rect 4028 19496 4034 19508
rect 4065 19499 4123 19505
rect 4065 19496 4077 19499
rect 4028 19468 4077 19496
rect 4028 19456 4034 19468
rect 4065 19465 4077 19468
rect 4111 19465 4123 19499
rect 4065 19459 4123 19465
rect 4982 19456 4988 19508
rect 5040 19456 5046 19508
rect 2774 19320 2780 19372
rect 2832 19360 2838 19372
rect 3142 19360 3148 19372
rect 2832 19332 3148 19360
rect 2832 19320 2838 19332
rect 3142 19320 3148 19332
rect 3200 19320 3206 19372
rect 4798 19320 4804 19372
rect 4856 19320 4862 19372
rect 2314 19252 2320 19304
rect 2372 19292 2378 19304
rect 3237 19295 3295 19301
rect 3237 19292 3249 19295
rect 2372 19264 3249 19292
rect 2372 19252 2378 19264
rect 3237 19261 3249 19264
rect 3283 19261 3295 19295
rect 3237 19255 3295 19261
rect 4338 19252 4344 19304
rect 4396 19292 4402 19304
rect 4617 19295 4675 19301
rect 4617 19292 4629 19295
rect 4396 19264 4629 19292
rect 4396 19252 4402 19264
rect 4617 19261 4629 19264
rect 4663 19261 4675 19295
rect 4617 19255 4675 19261
rect 1104 19066 5428 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 5428 19066
rect 1104 18992 5428 19014
rect 2314 18912 2320 18964
rect 2372 18912 2378 18964
rect 1670 18708 1676 18760
rect 1728 18748 1734 18760
rect 1949 18751 2007 18757
rect 1949 18748 1961 18751
rect 1728 18720 1961 18748
rect 1728 18708 1734 18720
rect 1949 18717 1961 18720
rect 1995 18717 2007 18751
rect 1949 18711 2007 18717
rect 2409 18751 2467 18757
rect 2409 18717 2421 18751
rect 2455 18748 2467 18751
rect 2774 18748 2780 18760
rect 2455 18720 2780 18748
rect 2455 18717 2467 18720
rect 2409 18711 2467 18717
rect 2774 18708 2780 18720
rect 2832 18708 2838 18760
rect 4706 18708 4712 18760
rect 4764 18708 4770 18760
rect 4062 18572 4068 18624
rect 4120 18572 4126 18624
rect 1104 18522 5428 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 5428 18522
rect 1104 18448 5428 18470
rect 2774 18368 2780 18420
rect 2832 18368 2838 18420
rect 4798 18408 4804 18420
rect 3804 18380 4804 18408
rect 3050 18340 3056 18352
rect 1412 18312 3056 18340
rect 1412 18281 1440 18312
rect 3050 18300 3056 18312
rect 3108 18340 3114 18352
rect 3108 18312 3740 18340
rect 3108 18300 3114 18312
rect 3712 18284 3740 18312
rect 1670 18281 1676 18284
rect 1397 18275 1455 18281
rect 1397 18241 1409 18275
rect 1443 18241 1455 18275
rect 1664 18272 1676 18281
rect 1631 18244 1676 18272
rect 1397 18235 1455 18241
rect 1664 18235 1676 18244
rect 1670 18232 1676 18235
rect 1728 18232 1734 18284
rect 3694 18232 3700 18284
rect 3752 18232 3758 18284
rect 3053 18207 3111 18213
rect 3053 18173 3065 18207
rect 3099 18204 3111 18207
rect 3804 18204 3832 18380
rect 4798 18368 4804 18380
rect 4856 18408 4862 18420
rect 5077 18411 5135 18417
rect 5077 18408 5089 18411
rect 4856 18380 5089 18408
rect 4856 18368 4862 18380
rect 5077 18377 5089 18380
rect 5123 18377 5135 18411
rect 5077 18371 5135 18377
rect 3964 18343 4022 18349
rect 3964 18309 3976 18343
rect 4010 18340 4022 18343
rect 4062 18340 4068 18352
rect 4010 18312 4068 18340
rect 4010 18309 4022 18312
rect 3964 18303 4022 18309
rect 4062 18300 4068 18312
rect 4120 18300 4126 18352
rect 3099 18176 3832 18204
rect 3099 18173 3111 18176
rect 3053 18167 3111 18173
rect 3605 18071 3663 18077
rect 3605 18037 3617 18071
rect 3651 18068 3663 18071
rect 4614 18068 4620 18080
rect 3651 18040 4620 18068
rect 3651 18037 3663 18040
rect 3605 18031 3663 18037
rect 4614 18028 4620 18040
rect 4672 18028 4678 18080
rect 1104 17978 5428 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 5428 17978
rect 1104 17904 5428 17926
rect 4157 17867 4215 17873
rect 4157 17833 4169 17867
rect 4203 17864 4215 17867
rect 4706 17864 4712 17876
rect 4203 17836 4712 17864
rect 4203 17833 4215 17836
rect 4157 17827 4215 17833
rect 4706 17824 4712 17836
rect 4764 17824 4770 17876
rect 1581 17799 1639 17805
rect 1581 17765 1593 17799
rect 1627 17796 1639 17799
rect 1670 17796 1676 17808
rect 1627 17768 1676 17796
rect 1627 17765 1639 17768
rect 1581 17759 1639 17765
rect 1670 17756 1676 17768
rect 1728 17796 1734 17808
rect 2685 17799 2743 17805
rect 1728 17768 2268 17796
rect 1728 17756 1734 17768
rect 658 17620 664 17672
rect 716 17660 722 17672
rect 2240 17669 2268 17768
rect 2685 17765 2697 17799
rect 2731 17796 2743 17799
rect 2731 17768 4752 17796
rect 2731 17765 2743 17768
rect 2685 17759 2743 17765
rect 4724 17740 4752 17768
rect 4614 17688 4620 17740
rect 4672 17688 4678 17740
rect 4706 17688 4712 17740
rect 4764 17728 4770 17740
rect 4801 17731 4859 17737
rect 4801 17728 4813 17731
rect 4764 17700 4813 17728
rect 4764 17688 4770 17700
rect 4801 17697 4813 17700
rect 4847 17728 4859 17731
rect 5258 17728 5264 17740
rect 4847 17700 5264 17728
rect 4847 17697 4859 17700
rect 4801 17691 4859 17697
rect 5258 17688 5264 17700
rect 5316 17688 5322 17740
rect 1397 17663 1455 17669
rect 1397 17660 1409 17663
rect 716 17632 1409 17660
rect 716 17620 722 17632
rect 1397 17629 1409 17632
rect 1443 17629 1455 17663
rect 1397 17623 1455 17629
rect 2225 17663 2283 17669
rect 2225 17629 2237 17663
rect 2271 17629 2283 17663
rect 2225 17623 2283 17629
rect 2774 17620 2780 17672
rect 2832 17660 2838 17672
rect 3145 17663 3203 17669
rect 3145 17660 3157 17663
rect 2832 17632 3157 17660
rect 2832 17620 2838 17632
rect 3145 17629 3157 17632
rect 3191 17629 3203 17663
rect 3145 17623 3203 17629
rect 4062 17484 4068 17536
rect 4120 17524 4126 17536
rect 4525 17527 4583 17533
rect 4525 17524 4537 17527
rect 4120 17496 4537 17524
rect 4120 17484 4126 17496
rect 4525 17493 4537 17496
rect 4571 17493 4583 17527
rect 4525 17487 4583 17493
rect 1104 17434 5428 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 5428 17434
rect 1104 17360 5428 17382
rect 3050 17144 3056 17196
rect 3108 17144 3114 17196
rect 3326 17193 3332 17196
rect 3320 17147 3332 17193
rect 3326 17144 3332 17147
rect 3384 17144 3390 17196
rect 4062 16940 4068 16992
rect 4120 16980 4126 16992
rect 4433 16983 4491 16989
rect 4433 16980 4445 16983
rect 4120 16952 4445 16980
rect 4120 16940 4126 16952
rect 4433 16949 4445 16952
rect 4479 16949 4491 16983
rect 4433 16943 4491 16949
rect 1104 16890 5428 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 5428 16890
rect 1104 16816 5428 16838
rect 2222 16736 2228 16788
rect 2280 16776 2286 16788
rect 2961 16779 3019 16785
rect 2961 16776 2973 16779
rect 2280 16748 2973 16776
rect 2280 16736 2286 16748
rect 2961 16745 2973 16748
rect 3007 16745 3019 16779
rect 2961 16739 3019 16745
rect 3326 16736 3332 16788
rect 3384 16736 3390 16788
rect 2869 16711 2927 16717
rect 2869 16677 2881 16711
rect 2915 16708 2927 16711
rect 2915 16680 3372 16708
rect 2915 16677 2927 16680
rect 2869 16671 2927 16677
rect 2130 16600 2136 16652
rect 2188 16640 2194 16652
rect 2314 16640 2320 16652
rect 2188 16612 2320 16640
rect 2188 16600 2194 16612
rect 2314 16600 2320 16612
rect 2372 16640 2378 16652
rect 2777 16643 2835 16649
rect 2777 16640 2789 16643
rect 2372 16612 2789 16640
rect 2372 16600 2378 16612
rect 2777 16609 2789 16612
rect 2823 16609 2835 16643
rect 2777 16603 2835 16609
rect 3053 16575 3111 16581
rect 3053 16541 3065 16575
rect 3099 16541 3111 16575
rect 3053 16535 3111 16541
rect 3068 16504 3096 16535
rect 3142 16532 3148 16584
rect 3200 16532 3206 16584
rect 3344 16581 3372 16680
rect 3878 16600 3884 16652
rect 3936 16640 3942 16652
rect 4062 16640 4068 16652
rect 3936 16612 4068 16640
rect 3936 16600 3942 16612
rect 4062 16600 4068 16612
rect 4120 16640 4126 16652
rect 4341 16643 4399 16649
rect 4341 16640 4353 16643
rect 4120 16612 4353 16640
rect 4120 16600 4126 16612
rect 4341 16609 4353 16612
rect 4387 16609 4399 16643
rect 4341 16603 4399 16609
rect 3329 16575 3387 16581
rect 3329 16541 3341 16575
rect 3375 16541 3387 16575
rect 3329 16535 3387 16541
rect 4798 16532 4804 16584
rect 4856 16532 4862 16584
rect 3789 16507 3847 16513
rect 3789 16504 3801 16507
rect 3068 16476 3801 16504
rect 3789 16473 3801 16476
rect 3835 16473 3847 16507
rect 3789 16467 3847 16473
rect 4985 16439 5043 16445
rect 4985 16405 4997 16439
rect 5031 16436 5043 16439
rect 5258 16436 5264 16448
rect 5031 16408 5264 16436
rect 5031 16405 5043 16408
rect 4985 16399 5043 16405
rect 5258 16396 5264 16408
rect 5316 16396 5322 16448
rect 1104 16346 5428 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 5428 16346
rect 1104 16272 5428 16294
rect 1946 16056 1952 16108
rect 2004 16096 2010 16108
rect 2041 16099 2099 16105
rect 2041 16096 2053 16099
rect 2004 16068 2053 16096
rect 2004 16056 2010 16068
rect 2041 16065 2053 16068
rect 2087 16065 2099 16099
rect 2041 16059 2099 16065
rect 2222 16056 2228 16108
rect 2280 16096 2286 16108
rect 2498 16096 2504 16108
rect 2280 16068 2504 16096
rect 2280 16056 2286 16068
rect 2498 16056 2504 16068
rect 2556 16056 2562 16108
rect 2038 15852 2044 15904
rect 2096 15852 2102 15904
rect 1104 15802 5428 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 5428 15802
rect 1104 15728 5428 15750
rect 2961 15691 3019 15697
rect 2961 15657 2973 15691
rect 3007 15688 3019 15691
rect 3142 15688 3148 15700
rect 3007 15660 3148 15688
rect 3007 15657 3019 15660
rect 2961 15651 3019 15657
rect 3142 15648 3148 15660
rect 3200 15648 3206 15700
rect 1397 15487 1455 15493
rect 1397 15453 1409 15487
rect 1443 15484 1455 15487
rect 3050 15484 3056 15496
rect 1443 15456 3056 15484
rect 1443 15453 1455 15456
rect 1397 15447 1455 15453
rect 3050 15444 3056 15456
rect 3108 15484 3114 15496
rect 3694 15484 3700 15496
rect 3108 15456 3700 15484
rect 3108 15444 3114 15456
rect 3694 15444 3700 15456
rect 3752 15444 3758 15496
rect 3970 15444 3976 15496
rect 4028 15484 4034 15496
rect 4617 15487 4675 15493
rect 4617 15484 4629 15487
rect 4028 15456 4629 15484
rect 4028 15444 4034 15456
rect 4617 15453 4629 15456
rect 4663 15453 4675 15487
rect 4617 15447 4675 15453
rect 1664 15419 1722 15425
rect 1664 15385 1676 15419
rect 1710 15416 1722 15419
rect 2038 15416 2044 15428
rect 1710 15388 2044 15416
rect 1710 15385 1722 15388
rect 1664 15379 1722 15385
rect 2038 15376 2044 15388
rect 2096 15376 2102 15428
rect 2590 15376 2596 15428
rect 2648 15416 2654 15428
rect 3145 15419 3203 15425
rect 3145 15416 3157 15419
rect 2648 15388 3157 15416
rect 2648 15376 2654 15388
rect 3145 15385 3157 15388
rect 3191 15385 3203 15419
rect 3145 15379 3203 15385
rect 3237 15419 3295 15425
rect 3237 15385 3249 15419
rect 3283 15416 3295 15419
rect 3283 15388 3464 15416
rect 3283 15385 3295 15388
rect 3237 15379 3295 15385
rect 2774 15308 2780 15360
rect 2832 15308 2838 15360
rect 3326 15308 3332 15360
rect 3384 15308 3390 15360
rect 3436 15348 3464 15388
rect 3510 15376 3516 15428
rect 3568 15376 3574 15428
rect 3878 15348 3884 15360
rect 3436 15320 3884 15348
rect 3878 15308 3884 15320
rect 3936 15308 3942 15360
rect 4062 15308 4068 15360
rect 4120 15308 4126 15360
rect 1104 15258 5428 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 5428 15258
rect 1104 15184 5428 15206
rect 1946 15104 1952 15156
rect 2004 15104 2010 15156
rect 2501 15147 2559 15153
rect 2501 15113 2513 15147
rect 2547 15144 2559 15147
rect 2866 15144 2872 15156
rect 2547 15116 2872 15144
rect 2547 15113 2559 15116
rect 2501 15107 2559 15113
rect 2866 15104 2872 15116
rect 2924 15144 2930 15156
rect 3510 15144 3516 15156
rect 2924 15116 3516 15144
rect 2924 15104 2930 15116
rect 3510 15104 3516 15116
rect 3568 15104 3574 15156
rect 2133 15079 2191 15085
rect 2133 15076 2145 15079
rect 1872 15048 2145 15076
rect 1872 15017 1900 15048
rect 2133 15045 2145 15048
rect 2179 15045 2191 15079
rect 2133 15039 2191 15045
rect 1857 15011 1915 15017
rect 1857 14977 1869 15011
rect 1903 14977 1915 15011
rect 1857 14971 1915 14977
rect 2038 14968 2044 15020
rect 2096 14968 2102 15020
rect 2317 15011 2375 15017
rect 2317 14977 2329 15011
rect 2363 14977 2375 15011
rect 2317 14971 2375 14977
rect 2332 14940 2360 14971
rect 2590 14968 2596 15020
rect 2648 14968 2654 15020
rect 2682 14968 2688 15020
rect 2740 14968 2746 15020
rect 2774 14940 2780 14952
rect 2332 14912 2780 14940
rect 2774 14900 2780 14912
rect 2832 14900 2838 14952
rect 3694 14764 3700 14816
rect 3752 14804 3758 14816
rect 3973 14807 4031 14813
rect 3973 14804 3985 14807
rect 3752 14776 3985 14804
rect 3752 14764 3758 14776
rect 3973 14773 3985 14776
rect 4019 14773 4031 14807
rect 3973 14767 4031 14773
rect 1104 14714 5428 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 5428 14714
rect 1104 14640 5428 14662
rect 2498 14560 2504 14612
rect 2556 14560 2562 14612
rect 2685 14603 2743 14609
rect 2685 14569 2697 14603
rect 2731 14569 2743 14603
rect 2685 14563 2743 14569
rect 2700 14532 2728 14563
rect 3970 14560 3976 14612
rect 4028 14600 4034 14612
rect 4065 14603 4123 14609
rect 4065 14600 4077 14603
rect 4028 14572 4077 14600
rect 4028 14560 4034 14572
rect 4065 14569 4077 14572
rect 4111 14569 4123 14603
rect 4065 14563 4123 14569
rect 2774 14532 2780 14544
rect 2700 14504 2780 14532
rect 2774 14492 2780 14504
rect 2832 14532 2838 14544
rect 3326 14532 3332 14544
rect 2832 14504 3332 14532
rect 2832 14492 2838 14504
rect 3326 14492 3332 14504
rect 3384 14532 3390 14544
rect 3384 14504 4476 14532
rect 3384 14492 3390 14504
rect 4448 14405 4476 14504
rect 4706 14424 4712 14476
rect 4764 14424 4770 14476
rect 3053 14399 3111 14405
rect 3053 14365 3065 14399
rect 3099 14365 3111 14399
rect 3053 14359 3111 14365
rect 4433 14399 4491 14405
rect 4433 14365 4445 14399
rect 4479 14365 4491 14399
rect 4433 14359 4491 14365
rect 2130 14288 2136 14340
rect 2188 14328 2194 14340
rect 2590 14328 2596 14340
rect 2188 14300 2596 14328
rect 2188 14288 2194 14300
rect 2590 14288 2596 14300
rect 2648 14337 2654 14340
rect 2648 14331 2711 14337
rect 2648 14297 2665 14331
rect 2699 14297 2711 14331
rect 2648 14291 2711 14297
rect 2648 14288 2654 14291
rect 2866 14288 2872 14340
rect 2924 14288 2930 14340
rect 3068 14260 3096 14359
rect 3605 14331 3663 14337
rect 3605 14297 3617 14331
rect 3651 14328 3663 14331
rect 4525 14331 4583 14337
rect 4525 14328 4537 14331
rect 3651 14300 4537 14328
rect 3651 14297 3663 14300
rect 3605 14291 3663 14297
rect 4525 14297 4537 14300
rect 4571 14297 4583 14331
rect 4525 14291 4583 14297
rect 4798 14260 4804 14272
rect 3068 14232 4804 14260
rect 4798 14220 4804 14232
rect 4856 14220 4862 14272
rect 1104 14170 5428 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 5428 14170
rect 1104 14096 5428 14118
rect 4798 14016 4804 14068
rect 4856 14056 4862 14068
rect 5077 14059 5135 14065
rect 5077 14056 5089 14059
rect 4856 14028 5089 14056
rect 4856 14016 4862 14028
rect 5077 14025 5089 14028
rect 5123 14025 5135 14059
rect 5077 14019 5135 14025
rect 3964 13991 4022 13997
rect 3964 13957 3976 13991
rect 4010 13988 4022 13991
rect 4062 13988 4068 14000
rect 4010 13960 4068 13988
rect 4010 13957 4022 13960
rect 3964 13951 4022 13957
rect 4062 13948 4068 13960
rect 4120 13948 4126 14000
rect 3050 13812 3056 13864
rect 3108 13852 3114 13864
rect 3694 13852 3700 13864
rect 3108 13824 3700 13852
rect 3108 13812 3114 13824
rect 3694 13812 3700 13824
rect 3752 13812 3758 13864
rect 1104 13626 5428 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 5428 13626
rect 1104 13552 5428 13574
rect 3789 13447 3847 13453
rect 3789 13413 3801 13447
rect 3835 13444 3847 13447
rect 4614 13444 4620 13456
rect 3835 13416 4620 13444
rect 3835 13413 3847 13416
rect 3789 13407 3847 13413
rect 4614 13404 4620 13416
rect 4672 13404 4678 13456
rect 4890 13404 4896 13456
rect 4948 13404 4954 13456
rect 2866 13336 2872 13388
rect 2924 13376 2930 13388
rect 3145 13379 3203 13385
rect 3145 13376 3157 13379
rect 2924 13348 3157 13376
rect 2924 13336 2930 13348
rect 3145 13345 3157 13348
rect 3191 13376 3203 13379
rect 4433 13379 4491 13385
rect 3191 13348 4200 13376
rect 3191 13345 3203 13348
rect 3145 13339 3203 13345
rect 4172 13317 4200 13348
rect 4433 13345 4445 13379
rect 4479 13376 4491 13379
rect 4706 13376 4712 13388
rect 4479 13348 4712 13376
rect 4479 13345 4491 13348
rect 4433 13339 4491 13345
rect 4706 13336 4712 13348
rect 4764 13336 4770 13388
rect 4157 13311 4215 13317
rect 4157 13277 4169 13311
rect 4203 13277 4215 13311
rect 4157 13271 4215 13277
rect 4798 13268 4804 13320
rect 4856 13308 4862 13320
rect 5077 13311 5135 13317
rect 5077 13308 5089 13311
rect 4856 13280 5089 13308
rect 4856 13268 4862 13280
rect 5077 13277 5089 13280
rect 5123 13277 5135 13311
rect 5077 13271 5135 13277
rect 2222 13132 2228 13184
rect 2280 13172 2286 13184
rect 2593 13175 2651 13181
rect 2593 13172 2605 13175
rect 2280 13144 2605 13172
rect 2280 13132 2286 13144
rect 2593 13141 2605 13144
rect 2639 13141 2651 13175
rect 2593 13135 2651 13141
rect 4249 13175 4307 13181
rect 4249 13141 4261 13175
rect 4295 13172 4307 13175
rect 4430 13172 4436 13184
rect 4295 13144 4436 13172
rect 4295 13141 4307 13144
rect 4249 13135 4307 13141
rect 4430 13132 4436 13144
rect 4488 13132 4494 13184
rect 1104 13082 5428 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 5428 13082
rect 1104 13008 5428 13030
rect 2222 12928 2228 12980
rect 2280 12928 2286 12980
rect 4430 12928 4436 12980
rect 4488 12928 4494 12980
rect 2409 12903 2467 12909
rect 2409 12869 2421 12903
rect 2455 12900 2467 12903
rect 2866 12900 2872 12912
rect 2455 12872 2872 12900
rect 2455 12869 2467 12872
rect 2409 12863 2467 12869
rect 2866 12860 2872 12872
rect 2924 12860 2930 12912
rect 2130 12792 2136 12844
rect 2188 12792 2194 12844
rect 2590 12792 2596 12844
rect 2648 12792 2654 12844
rect 4798 12724 4804 12776
rect 4856 12764 4862 12776
rect 4985 12767 5043 12773
rect 4985 12764 4997 12767
rect 4856 12736 4997 12764
rect 4856 12724 4862 12736
rect 4985 12733 4997 12736
rect 5031 12733 5043 12767
rect 4985 12727 5043 12733
rect 2406 12588 2412 12640
rect 2464 12588 2470 12640
rect 2682 12588 2688 12640
rect 2740 12628 2746 12640
rect 3881 12631 3939 12637
rect 3881 12628 3893 12631
rect 2740 12600 3893 12628
rect 2740 12588 2746 12600
rect 3881 12597 3893 12600
rect 3927 12597 3939 12631
rect 3881 12591 3939 12597
rect 1104 12538 5428 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 5428 12538
rect 1104 12464 5428 12486
rect 2866 12384 2872 12436
rect 2924 12424 2930 12436
rect 3053 12427 3111 12433
rect 3053 12424 3065 12427
rect 2924 12396 3065 12424
rect 2924 12384 2930 12396
rect 3053 12393 3065 12396
rect 3099 12393 3111 12427
rect 3053 12387 3111 12393
rect 2866 12248 2872 12300
rect 2924 12288 2930 12300
rect 2961 12291 3019 12297
rect 2961 12288 2973 12291
rect 2924 12260 2973 12288
rect 2924 12248 2930 12260
rect 2961 12257 2973 12260
rect 3007 12257 3019 12291
rect 2961 12251 3019 12257
rect 4525 12291 4583 12297
rect 4525 12257 4537 12291
rect 4571 12288 4583 12291
rect 4614 12288 4620 12300
rect 4571 12260 4620 12288
rect 4571 12257 4583 12260
rect 4525 12251 4583 12257
rect 4614 12248 4620 12260
rect 4672 12248 4678 12300
rect 1489 12223 1547 12229
rect 1489 12189 1501 12223
rect 1535 12220 1547 12223
rect 3050 12220 3056 12232
rect 1535 12192 3056 12220
rect 1535 12189 1547 12192
rect 1489 12183 1547 12189
rect 3050 12180 3056 12192
rect 3108 12180 3114 12232
rect 3142 12180 3148 12232
rect 3200 12180 3206 12232
rect 3237 12223 3295 12229
rect 3237 12189 3249 12223
rect 3283 12189 3295 12223
rect 3237 12183 3295 12189
rect 1756 12155 1814 12161
rect 1756 12121 1768 12155
rect 1802 12152 1814 12155
rect 2406 12152 2412 12164
rect 1802 12124 2412 12152
rect 1802 12121 1814 12124
rect 1756 12115 1814 12121
rect 2406 12112 2412 12124
rect 2464 12112 2470 12164
rect 2869 12087 2927 12093
rect 2869 12053 2881 12087
rect 2915 12084 2927 12087
rect 2958 12084 2964 12096
rect 2915 12056 2964 12084
rect 2915 12053 2927 12056
rect 2869 12047 2927 12053
rect 2958 12044 2964 12056
rect 3016 12084 3022 12096
rect 3252 12084 3280 12183
rect 3016 12056 3280 12084
rect 3016 12044 3022 12056
rect 3878 12044 3884 12096
rect 3936 12044 3942 12096
rect 1104 11994 5428 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 5428 11994
rect 1104 11920 5428 11942
rect 2038 11840 2044 11892
rect 2096 11880 2102 11892
rect 2866 11880 2872 11892
rect 2096 11852 2872 11880
rect 2096 11840 2102 11852
rect 1578 11772 1584 11824
rect 1636 11812 1642 11824
rect 2424 11821 2452 11852
rect 2866 11840 2872 11852
rect 2924 11880 2930 11892
rect 3234 11880 3240 11892
rect 2924 11852 3240 11880
rect 2924 11840 2930 11852
rect 3234 11840 3240 11852
rect 3292 11840 3298 11892
rect 4798 11840 4804 11892
rect 4856 11880 4862 11892
rect 4985 11883 5043 11889
rect 4985 11880 4997 11883
rect 4856 11852 4997 11880
rect 4856 11840 4862 11852
rect 4985 11849 4997 11852
rect 5031 11849 5043 11883
rect 4985 11843 5043 11849
rect 3878 11821 3884 11824
rect 2193 11815 2251 11821
rect 2193 11812 2205 11815
rect 1636 11784 2205 11812
rect 1636 11772 1642 11784
rect 2193 11781 2205 11784
rect 2239 11781 2251 11815
rect 2193 11775 2251 11781
rect 2409 11815 2467 11821
rect 2409 11781 2421 11815
rect 2455 11781 2467 11815
rect 3872 11812 3884 11821
rect 3839 11784 3884 11812
rect 2409 11775 2467 11781
rect 3872 11775 3884 11784
rect 3878 11772 3884 11775
rect 3936 11772 3942 11824
rect 3050 11704 3056 11756
rect 3108 11744 3114 11756
rect 3605 11747 3663 11753
rect 3605 11744 3617 11747
rect 3108 11716 3617 11744
rect 3108 11704 3114 11716
rect 3605 11713 3617 11716
rect 3651 11713 3663 11747
rect 3605 11707 3663 11713
rect 2038 11500 2044 11552
rect 2096 11500 2102 11552
rect 2222 11500 2228 11552
rect 2280 11500 2286 11552
rect 1104 11450 5428 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 5428 11450
rect 1104 11376 5428 11398
rect 1578 11296 1584 11348
rect 1636 11296 1642 11348
rect 4157 11271 4215 11277
rect 4157 11237 4169 11271
rect 4203 11268 4215 11271
rect 5350 11268 5356 11280
rect 4203 11240 5356 11268
rect 4203 11237 4215 11240
rect 4157 11231 4215 11237
rect 5350 11228 5356 11240
rect 5408 11228 5414 11280
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11101 1731 11135
rect 1673 11095 1731 11101
rect 1688 11064 1716 11095
rect 1762 11092 1768 11144
rect 1820 11092 1826 11144
rect 2038 11141 2044 11144
rect 2032 11132 2044 11141
rect 1999 11104 2044 11132
rect 2032 11095 2044 11104
rect 2038 11092 2044 11095
rect 2096 11092 2102 11144
rect 3142 11092 3148 11144
rect 3200 11092 3206 11144
rect 4341 11135 4399 11141
rect 4341 11101 4353 11135
rect 4387 11132 4399 11135
rect 5077 11135 5135 11141
rect 5077 11132 5089 11135
rect 4387 11104 5089 11132
rect 4387 11101 4399 11104
rect 4341 11095 4399 11101
rect 5077 11101 5089 11104
rect 5123 11132 5135 11135
rect 5258 11132 5264 11144
rect 5123 11104 5264 11132
rect 5123 11101 5135 11104
rect 5077 11095 5135 11101
rect 5258 11092 5264 11104
rect 5316 11092 5322 11144
rect 2130 11064 2136 11076
rect 1688 11036 2136 11064
rect 2130 11024 2136 11036
rect 2188 11064 2194 11076
rect 3160 11064 3188 11092
rect 2188 11036 3188 11064
rect 2188 11024 2194 11036
rect 2774 10956 2780 11008
rect 2832 10996 2838 11008
rect 3145 10999 3203 11005
rect 3145 10996 3157 10999
rect 2832 10968 3157 10996
rect 2832 10956 2838 10968
rect 3145 10965 3157 10968
rect 3191 10965 3203 10999
rect 3145 10959 3203 10965
rect 4433 10999 4491 11005
rect 4433 10965 4445 10999
rect 4479 10996 4491 10999
rect 4614 10996 4620 11008
rect 4479 10968 4620 10996
rect 4479 10965 4491 10968
rect 4433 10959 4491 10965
rect 4614 10956 4620 10968
rect 4672 10956 4678 11008
rect 1104 10906 5428 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 5428 10906
rect 1104 10832 5428 10854
rect 2222 10752 2228 10804
rect 2280 10792 2286 10804
rect 2317 10795 2375 10801
rect 2317 10792 2329 10795
rect 2280 10764 2329 10792
rect 2280 10752 2286 10764
rect 2317 10761 2329 10764
rect 2363 10761 2375 10795
rect 5077 10795 5135 10801
rect 2317 10755 2375 10761
rect 2516 10764 3556 10792
rect 1762 10684 1768 10736
rect 1820 10724 1826 10736
rect 2516 10724 2544 10764
rect 3418 10724 3424 10736
rect 1820 10696 2544 10724
rect 2608 10696 3424 10724
rect 1820 10684 1826 10696
rect 2406 10548 2412 10600
rect 2464 10588 2470 10600
rect 2608 10597 2636 10696
rect 3418 10684 3424 10696
rect 3476 10684 3482 10736
rect 3528 10656 3556 10764
rect 5077 10761 5089 10795
rect 5123 10792 5135 10795
rect 5258 10792 5264 10804
rect 5123 10764 5264 10792
rect 5123 10761 5135 10764
rect 5077 10755 5135 10761
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 3605 10727 3663 10733
rect 3605 10693 3617 10727
rect 3651 10724 3663 10727
rect 3942 10727 4000 10733
rect 3942 10724 3954 10727
rect 3651 10696 3954 10724
rect 3651 10693 3663 10696
rect 3605 10687 3663 10693
rect 3942 10693 3954 10696
rect 3988 10693 4000 10727
rect 3942 10687 4000 10693
rect 3697 10659 3755 10665
rect 3697 10656 3709 10659
rect 3528 10628 3709 10656
rect 3697 10625 3709 10628
rect 3743 10625 3755 10659
rect 3697 10619 3755 10625
rect 2501 10591 2559 10597
rect 2501 10588 2513 10591
rect 2464 10560 2513 10588
rect 2464 10548 2470 10560
rect 2501 10557 2513 10560
rect 2547 10557 2559 10591
rect 2501 10551 2559 10557
rect 2593 10591 2651 10597
rect 2593 10557 2605 10591
rect 2639 10557 2651 10591
rect 2593 10551 2651 10557
rect 2685 10591 2743 10597
rect 2685 10557 2697 10591
rect 2731 10557 2743 10591
rect 2685 10551 2743 10557
rect 2700 10452 2728 10551
rect 2774 10548 2780 10600
rect 2832 10548 2838 10600
rect 3050 10548 3056 10600
rect 3108 10548 3114 10600
rect 2958 10452 2964 10464
rect 2700 10424 2964 10452
rect 2958 10412 2964 10424
rect 3016 10412 3022 10464
rect 1104 10362 5428 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 5428 10362
rect 1104 10288 5428 10310
rect 3050 10208 3056 10260
rect 3108 10248 3114 10260
rect 4065 10251 4123 10257
rect 4065 10248 4077 10251
rect 3108 10220 4077 10248
rect 3108 10208 3114 10220
rect 4065 10217 4077 10220
rect 4111 10217 4123 10251
rect 4065 10211 4123 10217
rect 3053 10115 3111 10121
rect 3053 10081 3065 10115
rect 3099 10112 3111 10115
rect 3142 10112 3148 10124
rect 3099 10084 3148 10112
rect 3099 10081 3111 10084
rect 3053 10075 3111 10081
rect 3142 10072 3148 10084
rect 3200 10072 3206 10124
rect 4706 10072 4712 10124
rect 4764 10072 4770 10124
rect 2774 10004 2780 10056
rect 2832 10044 2838 10056
rect 3237 10047 3295 10053
rect 3237 10044 3249 10047
rect 2832 10016 3249 10044
rect 2832 10004 2838 10016
rect 3237 10013 3249 10016
rect 3283 10044 3295 10047
rect 4433 10047 4491 10053
rect 4433 10044 4445 10047
rect 3283 10016 4445 10044
rect 3283 10013 3295 10016
rect 3237 10007 3295 10013
rect 4433 10013 4445 10016
rect 4479 10013 4491 10047
rect 4433 10007 4491 10013
rect 1394 9936 1400 9988
rect 1452 9976 1458 9988
rect 1762 9976 1768 9988
rect 1452 9948 1768 9976
rect 1452 9936 1458 9948
rect 1762 9936 1768 9948
rect 1820 9976 1826 9988
rect 2498 9976 2504 9988
rect 1820 9948 2504 9976
rect 1820 9936 1826 9948
rect 2498 9936 2504 9948
rect 2556 9936 2562 9988
rect 2958 9936 2964 9988
rect 3016 9976 3022 9988
rect 3605 9979 3663 9985
rect 3605 9976 3617 9979
rect 3016 9948 3617 9976
rect 3016 9936 3022 9948
rect 3605 9945 3617 9948
rect 3651 9945 3663 9979
rect 3605 9939 3663 9945
rect 4525 9979 4583 9985
rect 4525 9945 4537 9979
rect 4571 9976 4583 9979
rect 4614 9976 4620 9988
rect 4571 9948 4620 9976
rect 4571 9945 4583 9948
rect 4525 9939 4583 9945
rect 4614 9936 4620 9948
rect 4672 9936 4678 9988
rect 3326 9868 3332 9920
rect 3384 9868 3390 9920
rect 3418 9868 3424 9920
rect 3476 9868 3482 9920
rect 1104 9818 5428 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 5428 9818
rect 1104 9744 5428 9766
rect 2498 9664 2504 9716
rect 2556 9704 2562 9716
rect 3973 9707 4031 9713
rect 3973 9704 3985 9707
rect 2556 9676 3985 9704
rect 2556 9664 2562 9676
rect 3973 9673 3985 9676
rect 4019 9673 4031 9707
rect 3973 9667 4031 9673
rect 2148 9608 2360 9636
rect 2148 9577 2176 9608
rect 2133 9571 2191 9577
rect 2133 9537 2145 9571
rect 2179 9537 2191 9571
rect 2133 9531 2191 9537
rect 2225 9571 2283 9577
rect 2225 9537 2237 9571
rect 2271 9537 2283 9571
rect 2225 9531 2283 9537
rect 2240 9432 2268 9531
rect 2332 9500 2360 9608
rect 2682 9596 2688 9648
rect 2740 9596 2746 9648
rect 2406 9528 2412 9580
rect 2464 9568 2470 9580
rect 3326 9568 3332 9580
rect 2464 9540 3332 9568
rect 2464 9528 2470 9540
rect 3326 9528 3332 9540
rect 3384 9528 3390 9580
rect 3418 9500 3424 9512
rect 2332 9472 3424 9500
rect 3418 9460 3424 9472
rect 3476 9460 3482 9512
rect 2958 9432 2964 9444
rect 2240 9404 2964 9432
rect 2958 9392 2964 9404
rect 3016 9392 3022 9444
rect 2593 9367 2651 9373
rect 2593 9333 2605 9367
rect 2639 9364 2651 9367
rect 3050 9364 3056 9376
rect 2639 9336 3056 9364
rect 2639 9333 2651 9336
rect 2593 9327 2651 9333
rect 3050 9324 3056 9336
rect 3108 9324 3114 9376
rect 1104 9274 5428 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 5428 9274
rect 1104 9200 5428 9222
rect 3050 9120 3056 9172
rect 3108 9120 3114 9172
rect 2777 9095 2835 9101
rect 2777 9061 2789 9095
rect 2823 9092 2835 9095
rect 3326 9092 3332 9104
rect 2823 9064 3332 9092
rect 2823 9061 2835 9064
rect 2777 9055 2835 9061
rect 3326 9052 3332 9064
rect 3384 9092 3390 9104
rect 3384 9064 3648 9092
rect 3384 9052 3390 9064
rect 1394 8916 1400 8968
rect 1452 8916 1458 8968
rect 2958 8916 2964 8968
rect 3016 8956 3022 8968
rect 3329 8959 3387 8965
rect 3329 8956 3341 8959
rect 3016 8928 3341 8956
rect 3016 8916 3022 8928
rect 3329 8925 3341 8928
rect 3375 8925 3387 8959
rect 3329 8919 3387 8925
rect 3620 8900 3648 9064
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8956 5135 8959
rect 5258 8956 5264 8968
rect 5123 8928 5264 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 5258 8916 5264 8928
rect 5316 8916 5322 8968
rect 1664 8891 1722 8897
rect 1664 8857 1676 8891
rect 1710 8888 1722 8891
rect 1710 8860 2912 8888
rect 1710 8857 1722 8860
rect 1664 8851 1722 8857
rect 2884 8829 2912 8860
rect 3234 8848 3240 8900
rect 3292 8848 3298 8900
rect 3418 8848 3424 8900
rect 3476 8848 3482 8900
rect 3602 8848 3608 8900
rect 3660 8848 3666 8900
rect 2869 8823 2927 8829
rect 2869 8789 2881 8823
rect 2915 8789 2927 8823
rect 2869 8783 2927 8789
rect 3037 8823 3095 8829
rect 3037 8789 3049 8823
rect 3083 8820 3095 8823
rect 3329 8823 3387 8829
rect 3329 8820 3341 8823
rect 3083 8792 3341 8820
rect 3083 8789 3095 8792
rect 3037 8783 3095 8789
rect 3329 8789 3341 8792
rect 3375 8789 3387 8823
rect 3329 8783 3387 8789
rect 4433 8823 4491 8829
rect 4433 8789 4445 8823
rect 4479 8820 4491 8823
rect 4614 8820 4620 8832
rect 4479 8792 4620 8820
rect 4479 8789 4491 8792
rect 4433 8783 4491 8789
rect 4614 8780 4620 8792
rect 4672 8780 4678 8832
rect 1104 8730 5428 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 5428 8730
rect 1104 8656 5428 8678
rect 5077 8619 5135 8625
rect 5077 8585 5089 8619
rect 5123 8616 5135 8619
rect 5258 8616 5264 8628
rect 5123 8588 5264 8616
rect 5123 8585 5135 8588
rect 5077 8579 5135 8585
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 3605 8551 3663 8557
rect 3605 8517 3617 8551
rect 3651 8548 3663 8551
rect 3942 8551 4000 8557
rect 3942 8548 3954 8551
rect 3651 8520 3954 8548
rect 3651 8517 3663 8520
rect 3605 8511 3663 8517
rect 3942 8517 3954 8520
rect 3988 8517 4000 8551
rect 3942 8511 4000 8517
rect 1394 8440 1400 8492
rect 1452 8480 1458 8492
rect 3697 8483 3755 8489
rect 3697 8480 3709 8483
rect 1452 8452 3709 8480
rect 1452 8440 1458 8452
rect 3697 8449 3709 8452
rect 3743 8449 3755 8483
rect 3697 8443 3755 8449
rect 3050 8372 3056 8424
rect 3108 8372 3114 8424
rect 1104 8186 5428 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 5428 8186
rect 1104 8112 5428 8134
rect 3050 8032 3056 8084
rect 3108 8072 3114 8084
rect 3973 8075 4031 8081
rect 3973 8072 3985 8075
rect 3108 8044 3985 8072
rect 3108 8032 3114 8044
rect 3973 8041 3985 8044
rect 4019 8041 4031 8075
rect 3973 8035 4031 8041
rect 4525 7939 4583 7945
rect 4525 7905 4537 7939
rect 4571 7936 4583 7939
rect 4706 7936 4712 7948
rect 4571 7908 4712 7936
rect 4571 7905 4583 7908
rect 4525 7899 4583 7905
rect 4706 7896 4712 7908
rect 4764 7896 4770 7948
rect 3602 7828 3608 7880
rect 3660 7868 3666 7880
rect 4341 7871 4399 7877
rect 4341 7868 4353 7871
rect 3660 7840 4353 7868
rect 3660 7828 3666 7840
rect 4341 7837 4353 7840
rect 4387 7837 4399 7871
rect 4341 7831 4399 7837
rect 4433 7871 4491 7877
rect 4433 7837 4445 7871
rect 4479 7868 4491 7871
rect 4614 7868 4620 7880
rect 4479 7840 4620 7868
rect 4479 7837 4491 7840
rect 4433 7831 4491 7837
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7868 4859 7871
rect 5258 7868 5264 7880
rect 4847 7840 5264 7868
rect 4847 7837 4859 7840
rect 4801 7831 4859 7837
rect 5258 7828 5264 7840
rect 5316 7828 5322 7880
rect 4985 7735 5043 7741
rect 4985 7701 4997 7735
rect 5031 7732 5043 7735
rect 5810 7732 5816 7744
rect 5031 7704 5816 7732
rect 5031 7701 5043 7704
rect 4985 7695 5043 7701
rect 5810 7692 5816 7704
rect 5868 7692 5874 7744
rect 1104 7642 5428 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 5428 7642
rect 1104 7568 5428 7590
rect 2958 7284 2964 7336
rect 3016 7324 3022 7336
rect 3053 7327 3111 7333
rect 3053 7324 3065 7327
rect 3016 7296 3065 7324
rect 3016 7284 3022 7296
rect 3053 7293 3065 7296
rect 3099 7293 3111 7327
rect 3053 7287 3111 7293
rect 3234 7216 3240 7268
rect 3292 7256 3298 7268
rect 3329 7259 3387 7265
rect 3329 7256 3341 7259
rect 3292 7228 3341 7256
rect 3292 7216 3298 7228
rect 3329 7225 3341 7228
rect 3375 7225 3387 7259
rect 3329 7219 3387 7225
rect 3510 7148 3516 7200
rect 3568 7148 3574 7200
rect 1104 7098 5428 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 5428 7098
rect 1104 7024 5428 7046
rect 1394 6808 1400 6860
rect 1452 6808 1458 6860
rect 3234 6808 3240 6860
rect 3292 6848 3298 6860
rect 3329 6851 3387 6857
rect 3329 6848 3341 6851
rect 3292 6820 3341 6848
rect 3292 6808 3298 6820
rect 3329 6817 3341 6820
rect 3375 6817 3387 6851
rect 3329 6811 3387 6817
rect 2869 6783 2927 6789
rect 2869 6780 2881 6783
rect 2792 6752 2881 6780
rect 1664 6715 1722 6721
rect 1664 6681 1676 6715
rect 1710 6712 1722 6715
rect 2038 6712 2044 6724
rect 1710 6684 2044 6712
rect 1710 6681 1722 6684
rect 1664 6675 1722 6681
rect 2038 6672 2044 6684
rect 2096 6672 2102 6724
rect 2792 6656 2820 6752
rect 2869 6749 2881 6752
rect 2915 6780 2927 6783
rect 3418 6780 3424 6792
rect 2915 6752 3424 6780
rect 2915 6749 2927 6752
rect 2869 6743 2927 6749
rect 3418 6740 3424 6752
rect 3476 6740 3482 6792
rect 2958 6672 2964 6724
rect 3016 6712 3022 6724
rect 4614 6712 4620 6724
rect 3016 6684 4620 6712
rect 3016 6672 3022 6684
rect 4614 6672 4620 6684
rect 4672 6672 4678 6724
rect 2774 6604 2780 6656
rect 2832 6604 2838 6656
rect 3050 6604 3056 6656
rect 3108 6604 3114 6656
rect 1104 6554 5428 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 5428 6554
rect 1104 6480 5428 6502
rect 2038 6400 2044 6452
rect 2096 6400 2102 6452
rect 1394 6332 1400 6384
rect 1452 6372 1458 6384
rect 2682 6372 2688 6384
rect 1452 6344 2688 6372
rect 1452 6332 1458 6344
rect 2682 6332 2688 6344
rect 2740 6372 2746 6384
rect 2740 6344 3464 6372
rect 2740 6332 2746 6344
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6304 2283 6307
rect 3050 6304 3056 6316
rect 2271 6276 3056 6304
rect 2271 6273 2283 6276
rect 2225 6267 2283 6273
rect 3050 6264 3056 6276
rect 3108 6264 3114 6316
rect 3436 6313 3464 6344
rect 3510 6332 3516 6384
rect 3568 6372 3574 6384
rect 3666 6375 3724 6381
rect 3666 6372 3678 6375
rect 3568 6344 3678 6372
rect 3568 6332 3574 6344
rect 3666 6341 3678 6344
rect 3712 6341 3724 6375
rect 3666 6335 3724 6341
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6273 3479 6307
rect 3421 6267 3479 6273
rect 2501 6239 2559 6245
rect 2501 6205 2513 6239
rect 2547 6236 2559 6239
rect 2958 6236 2964 6248
rect 2547 6208 2964 6236
rect 2547 6205 2559 6208
rect 2501 6199 2559 6205
rect 2958 6196 2964 6208
rect 3016 6196 3022 6248
rect 2409 6171 2467 6177
rect 2409 6137 2421 6171
rect 2455 6168 2467 6171
rect 2774 6168 2780 6180
rect 2455 6140 2780 6168
rect 2455 6137 2467 6140
rect 2409 6131 2467 6137
rect 2774 6128 2780 6140
rect 2832 6128 2838 6180
rect 4614 6060 4620 6112
rect 4672 6100 4678 6112
rect 4801 6103 4859 6109
rect 4801 6100 4813 6103
rect 4672 6072 4813 6100
rect 4672 6060 4678 6072
rect 4801 6069 4813 6072
rect 4847 6069 4859 6103
rect 4801 6063 4859 6069
rect 1104 6010 5428 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 5428 6010
rect 1104 5936 5428 5958
rect 3602 5652 3608 5704
rect 3660 5652 3666 5704
rect 5077 5695 5135 5701
rect 5077 5661 5089 5695
rect 5123 5692 5135 5695
rect 5350 5692 5356 5704
rect 5123 5664 5356 5692
rect 5123 5661 5135 5664
rect 5077 5655 5135 5661
rect 5350 5652 5356 5664
rect 5408 5652 5414 5704
rect 2958 5516 2964 5568
rect 3016 5516 3022 5568
rect 4433 5559 4491 5565
rect 4433 5525 4445 5559
rect 4479 5556 4491 5559
rect 4706 5556 4712 5568
rect 4479 5528 4712 5556
rect 4479 5525 4491 5528
rect 4433 5519 4491 5525
rect 4706 5516 4712 5528
rect 4764 5516 4770 5568
rect 1104 5466 5428 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 5428 5466
rect 1104 5392 5428 5414
rect 2958 5312 2964 5364
rect 3016 5352 3022 5364
rect 3237 5355 3295 5361
rect 3237 5352 3249 5355
rect 3016 5324 3249 5352
rect 3016 5312 3022 5324
rect 3237 5321 3249 5324
rect 3283 5321 3295 5355
rect 3237 5315 3295 5321
rect 2682 5244 2688 5296
rect 2740 5284 2746 5296
rect 2740 5256 3740 5284
rect 2740 5244 2746 5256
rect 2774 5176 2780 5228
rect 2832 5216 2838 5228
rect 3712 5225 3740 5256
rect 3970 5225 3976 5228
rect 3145 5219 3203 5225
rect 3145 5216 3157 5219
rect 2832 5188 3157 5216
rect 2832 5176 2838 5188
rect 3145 5185 3157 5188
rect 3191 5185 3203 5219
rect 3145 5179 3203 5185
rect 3697 5219 3755 5225
rect 3697 5185 3709 5219
rect 3743 5185 3755 5219
rect 3697 5179 3755 5185
rect 3964 5179 3976 5225
rect 3970 5176 3976 5179
rect 4028 5176 4034 5228
rect 3421 5151 3479 5157
rect 3421 5117 3433 5151
rect 3467 5117 3479 5151
rect 3421 5111 3479 5117
rect 2498 4972 2504 5024
rect 2556 5012 2562 5024
rect 2777 5015 2835 5021
rect 2777 5012 2789 5015
rect 2556 4984 2789 5012
rect 2556 4972 2562 4984
rect 2777 4981 2789 4984
rect 2823 4981 2835 5015
rect 3436 5012 3464 5111
rect 4798 5012 4804 5024
rect 3436 4984 4804 5012
rect 2777 4975 2835 4981
rect 4798 4972 4804 4984
rect 4856 4972 4862 5024
rect 5077 5015 5135 5021
rect 5077 4981 5089 5015
rect 5123 5012 5135 5015
rect 5350 5012 5356 5024
rect 5123 4984 5356 5012
rect 5123 4981 5135 4984
rect 5077 4975 5135 4981
rect 5350 4972 5356 4984
rect 5408 4972 5414 5024
rect 1104 4922 5428 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 5428 4922
rect 1104 4848 5428 4870
rect 3970 4768 3976 4820
rect 4028 4808 4034 4820
rect 4249 4811 4307 4817
rect 4249 4808 4261 4811
rect 4028 4780 4261 4808
rect 4028 4768 4034 4780
rect 4249 4777 4261 4780
rect 4295 4777 4307 4811
rect 4249 4771 4307 4777
rect 4706 4632 4712 4684
rect 4764 4632 4770 4684
rect 4798 4632 4804 4684
rect 4856 4632 4862 4684
rect 2225 4607 2283 4613
rect 2225 4573 2237 4607
rect 2271 4604 2283 4607
rect 2271 4576 2728 4604
rect 2271 4573 2283 4576
rect 2225 4567 2283 4573
rect 2700 4548 2728 4576
rect 4614 4564 4620 4616
rect 4672 4564 4678 4616
rect 2498 4545 2504 4548
rect 2492 4536 2504 4545
rect 2459 4508 2504 4536
rect 2492 4499 2504 4508
rect 2498 4496 2504 4499
rect 2556 4496 2562 4548
rect 2682 4496 2688 4548
rect 2740 4496 2746 4548
rect 3602 4428 3608 4480
rect 3660 4468 3666 4480
rect 4154 4468 4160 4480
rect 3660 4440 4160 4468
rect 3660 4428 3666 4440
rect 4154 4428 4160 4440
rect 4212 4428 4218 4480
rect 1104 4378 5428 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 5428 4378
rect 1104 4304 5428 4326
rect 4154 4088 4160 4140
rect 4212 4128 4218 4140
rect 4801 4131 4859 4137
rect 4801 4128 4813 4131
rect 4212 4100 4813 4128
rect 4212 4088 4218 4100
rect 4801 4097 4813 4100
rect 4847 4097 4859 4131
rect 4801 4091 4859 4097
rect 4985 3995 5043 4001
rect 4985 3961 4997 3995
rect 5031 3992 5043 3995
rect 5258 3992 5264 4004
rect 5031 3964 5264 3992
rect 5031 3961 5043 3964
rect 4985 3955 5043 3961
rect 5258 3952 5264 3964
rect 5316 3952 5322 4004
rect 1104 3834 5428 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 5428 3834
rect 1104 3760 5428 3782
rect 1104 3290 5428 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 5428 3290
rect 1104 3216 5428 3238
rect 1104 2746 5428 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 5428 2746
rect 1104 2672 5428 2694
rect 5077 2431 5135 2437
rect 5077 2397 5089 2431
rect 5123 2428 5135 2431
rect 5350 2428 5356 2440
rect 5123 2400 5356 2428
rect 5123 2397 5135 2400
rect 5077 2391 5135 2397
rect 5350 2388 5356 2400
rect 5408 2388 5414 2440
rect 4893 2295 4951 2301
rect 4893 2261 4905 2295
rect 4939 2292 4951 2295
rect 6362 2292 6368 2304
rect 4939 2264 6368 2292
rect 4939 2261 4951 2264
rect 4893 2255 4951 2261
rect 6362 2252 6368 2264
rect 6420 2252 6426 2304
rect 1104 2202 5428 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 5428 2202
rect 1104 2128 5428 2150
<< via1 >>
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 5264 21632 5316 21684
rect 4804 21539 4856 21548
rect 4804 21505 4813 21539
rect 4813 21505 4847 21539
rect 4847 21505 4856 21539
rect 4804 21496 4856 21505
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 4804 20952 4856 21004
rect 4620 20748 4672 20800
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 4804 20544 4856 20596
rect 2504 20451 2556 20460
rect 2504 20417 2538 20451
rect 2538 20417 2556 20451
rect 2504 20408 2556 20417
rect 3700 20451 3752 20460
rect 3700 20417 3709 20451
rect 3709 20417 3743 20451
rect 3743 20417 3752 20451
rect 3700 20408 3752 20417
rect 3976 20451 4028 20460
rect 3976 20417 4010 20451
rect 4010 20417 4028 20451
rect 3976 20408 4028 20417
rect 3608 20247 3660 20256
rect 3608 20213 3617 20247
rect 3617 20213 3651 20247
rect 3651 20213 3660 20247
rect 3608 20204 3660 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 2504 20000 2556 20052
rect 3608 19907 3660 19916
rect 3608 19873 3617 19907
rect 3617 19873 3651 19907
rect 3651 19873 3660 19907
rect 3608 19864 3660 19873
rect 2780 19839 2832 19848
rect 2780 19805 2789 19839
rect 2789 19805 2823 19839
rect 2823 19805 2832 19839
rect 2780 19796 2832 19805
rect 2872 19839 2924 19848
rect 2872 19805 2881 19839
rect 2881 19805 2915 19839
rect 2915 19805 2924 19839
rect 5264 19864 5316 19916
rect 2872 19796 2924 19805
rect 4620 19728 4672 19780
rect 2964 19660 3016 19712
rect 4344 19660 4396 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 2872 19499 2924 19508
rect 2872 19465 2881 19499
rect 2881 19465 2915 19499
rect 2915 19465 2924 19499
rect 2872 19456 2924 19465
rect 2964 19499 3016 19508
rect 2964 19465 2973 19499
rect 2973 19465 3007 19499
rect 3007 19465 3016 19499
rect 2964 19456 3016 19465
rect 3976 19456 4028 19508
rect 4988 19499 5040 19508
rect 4988 19465 4997 19499
rect 4997 19465 5031 19499
rect 5031 19465 5040 19499
rect 4988 19456 5040 19465
rect 2780 19363 2832 19372
rect 2780 19329 2789 19363
rect 2789 19329 2823 19363
rect 2823 19329 2832 19363
rect 2780 19320 2832 19329
rect 3148 19320 3200 19372
rect 4804 19363 4856 19372
rect 4804 19329 4813 19363
rect 4813 19329 4847 19363
rect 4847 19329 4856 19363
rect 4804 19320 4856 19329
rect 2320 19252 2372 19304
rect 4344 19252 4396 19304
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 2320 18955 2372 18964
rect 2320 18921 2329 18955
rect 2329 18921 2363 18955
rect 2363 18921 2372 18955
rect 2320 18912 2372 18921
rect 1676 18708 1728 18760
rect 2780 18708 2832 18760
rect 4712 18751 4764 18760
rect 4712 18717 4721 18751
rect 4721 18717 4755 18751
rect 4755 18717 4764 18751
rect 4712 18708 4764 18717
rect 4068 18615 4120 18624
rect 4068 18581 4077 18615
rect 4077 18581 4111 18615
rect 4111 18581 4120 18615
rect 4068 18572 4120 18581
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 2780 18411 2832 18420
rect 2780 18377 2789 18411
rect 2789 18377 2823 18411
rect 2823 18377 2832 18411
rect 2780 18368 2832 18377
rect 3056 18300 3108 18352
rect 1676 18275 1728 18284
rect 1676 18241 1710 18275
rect 1710 18241 1728 18275
rect 1676 18232 1728 18241
rect 3700 18275 3752 18284
rect 3700 18241 3709 18275
rect 3709 18241 3743 18275
rect 3743 18241 3752 18275
rect 3700 18232 3752 18241
rect 4804 18368 4856 18420
rect 4068 18300 4120 18352
rect 4620 18028 4672 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 4712 17824 4764 17876
rect 1676 17756 1728 17808
rect 664 17620 716 17672
rect 4620 17731 4672 17740
rect 4620 17697 4629 17731
rect 4629 17697 4663 17731
rect 4663 17697 4672 17731
rect 4620 17688 4672 17697
rect 4712 17688 4764 17740
rect 5264 17688 5316 17740
rect 2780 17620 2832 17672
rect 4068 17484 4120 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 3056 17187 3108 17196
rect 3056 17153 3065 17187
rect 3065 17153 3099 17187
rect 3099 17153 3108 17187
rect 3056 17144 3108 17153
rect 3332 17187 3384 17196
rect 3332 17153 3366 17187
rect 3366 17153 3384 17187
rect 3332 17144 3384 17153
rect 4068 16940 4120 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 2228 16736 2280 16788
rect 3332 16779 3384 16788
rect 3332 16745 3341 16779
rect 3341 16745 3375 16779
rect 3375 16745 3384 16779
rect 3332 16736 3384 16745
rect 2136 16600 2188 16652
rect 2320 16600 2372 16652
rect 3148 16575 3200 16584
rect 3148 16541 3157 16575
rect 3157 16541 3191 16575
rect 3191 16541 3200 16575
rect 3148 16532 3200 16541
rect 3884 16600 3936 16652
rect 4068 16600 4120 16652
rect 4804 16575 4856 16584
rect 4804 16541 4813 16575
rect 4813 16541 4847 16575
rect 4847 16541 4856 16575
rect 4804 16532 4856 16541
rect 5264 16396 5316 16448
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 1952 16056 2004 16108
rect 2228 16099 2280 16108
rect 2228 16065 2237 16099
rect 2237 16065 2271 16099
rect 2271 16065 2280 16099
rect 2228 16056 2280 16065
rect 2504 16056 2556 16108
rect 2044 15895 2096 15904
rect 2044 15861 2053 15895
rect 2053 15861 2087 15895
rect 2087 15861 2096 15895
rect 2044 15852 2096 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 3148 15648 3200 15700
rect 3056 15444 3108 15496
rect 3700 15444 3752 15496
rect 3976 15444 4028 15496
rect 2044 15376 2096 15428
rect 2596 15376 2648 15428
rect 2780 15351 2832 15360
rect 2780 15317 2789 15351
rect 2789 15317 2823 15351
rect 2823 15317 2832 15351
rect 2780 15308 2832 15317
rect 3332 15351 3384 15360
rect 3332 15317 3341 15351
rect 3341 15317 3375 15351
rect 3375 15317 3384 15351
rect 3332 15308 3384 15317
rect 3516 15419 3568 15428
rect 3516 15385 3525 15419
rect 3525 15385 3559 15419
rect 3559 15385 3568 15419
rect 3516 15376 3568 15385
rect 3884 15308 3936 15360
rect 4068 15351 4120 15360
rect 4068 15317 4077 15351
rect 4077 15317 4111 15351
rect 4111 15317 4120 15351
rect 4068 15308 4120 15317
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 1952 15147 2004 15156
rect 1952 15113 1961 15147
rect 1961 15113 1995 15147
rect 1995 15113 2004 15147
rect 1952 15104 2004 15113
rect 2872 15104 2924 15156
rect 3516 15104 3568 15156
rect 2044 15011 2096 15020
rect 2044 14977 2053 15011
rect 2053 14977 2087 15011
rect 2087 14977 2096 15011
rect 2044 14968 2096 14977
rect 2596 15011 2648 15020
rect 2596 14977 2605 15011
rect 2605 14977 2639 15011
rect 2639 14977 2648 15011
rect 2596 14968 2648 14977
rect 2688 15011 2740 15020
rect 2688 14977 2697 15011
rect 2697 14977 2731 15011
rect 2731 14977 2740 15011
rect 2688 14968 2740 14977
rect 2780 14900 2832 14952
rect 3700 14764 3752 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 2504 14603 2556 14612
rect 2504 14569 2513 14603
rect 2513 14569 2547 14603
rect 2547 14569 2556 14603
rect 2504 14560 2556 14569
rect 3976 14560 4028 14612
rect 2780 14492 2832 14544
rect 3332 14492 3384 14544
rect 4712 14467 4764 14476
rect 4712 14433 4721 14467
rect 4721 14433 4755 14467
rect 4755 14433 4764 14467
rect 4712 14424 4764 14433
rect 2136 14288 2188 14340
rect 2596 14288 2648 14340
rect 2872 14331 2924 14340
rect 2872 14297 2881 14331
rect 2881 14297 2915 14331
rect 2915 14297 2924 14331
rect 2872 14288 2924 14297
rect 4804 14220 4856 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 4804 14016 4856 14068
rect 4068 13948 4120 14000
rect 3056 13812 3108 13864
rect 3700 13855 3752 13864
rect 3700 13821 3709 13855
rect 3709 13821 3743 13855
rect 3743 13821 3752 13855
rect 3700 13812 3752 13821
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 4620 13404 4672 13456
rect 4896 13447 4948 13456
rect 4896 13413 4905 13447
rect 4905 13413 4939 13447
rect 4939 13413 4948 13447
rect 4896 13404 4948 13413
rect 2872 13336 2924 13388
rect 4712 13336 4764 13388
rect 4804 13268 4856 13320
rect 2228 13132 2280 13184
rect 4436 13132 4488 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 2228 12971 2280 12980
rect 2228 12937 2237 12971
rect 2237 12937 2271 12971
rect 2271 12937 2280 12971
rect 2228 12928 2280 12937
rect 4436 12971 4488 12980
rect 4436 12937 4445 12971
rect 4445 12937 4479 12971
rect 4479 12937 4488 12971
rect 4436 12928 4488 12937
rect 2872 12860 2924 12912
rect 2136 12835 2188 12844
rect 2136 12801 2145 12835
rect 2145 12801 2179 12835
rect 2179 12801 2188 12835
rect 2136 12792 2188 12801
rect 2596 12835 2648 12844
rect 2596 12801 2605 12835
rect 2605 12801 2639 12835
rect 2639 12801 2648 12835
rect 2596 12792 2648 12801
rect 4804 12724 4856 12776
rect 2412 12631 2464 12640
rect 2412 12597 2421 12631
rect 2421 12597 2455 12631
rect 2455 12597 2464 12631
rect 2412 12588 2464 12597
rect 2688 12588 2740 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 2872 12384 2924 12436
rect 2872 12248 2924 12300
rect 4620 12248 4672 12300
rect 3056 12180 3108 12232
rect 3148 12223 3200 12232
rect 3148 12189 3157 12223
rect 3157 12189 3191 12223
rect 3191 12189 3200 12223
rect 3148 12180 3200 12189
rect 2412 12112 2464 12164
rect 2964 12044 3016 12096
rect 3884 12087 3936 12096
rect 3884 12053 3893 12087
rect 3893 12053 3927 12087
rect 3927 12053 3936 12087
rect 3884 12044 3936 12053
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 2044 11840 2096 11892
rect 1584 11772 1636 11824
rect 2872 11840 2924 11892
rect 3240 11840 3292 11892
rect 4804 11840 4856 11892
rect 3884 11815 3936 11824
rect 3884 11781 3918 11815
rect 3918 11781 3936 11815
rect 3884 11772 3936 11781
rect 3056 11704 3108 11756
rect 2044 11543 2096 11552
rect 2044 11509 2053 11543
rect 2053 11509 2087 11543
rect 2087 11509 2096 11543
rect 2044 11500 2096 11509
rect 2228 11543 2280 11552
rect 2228 11509 2237 11543
rect 2237 11509 2271 11543
rect 2271 11509 2280 11543
rect 2228 11500 2280 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 1584 11339 1636 11348
rect 1584 11305 1593 11339
rect 1593 11305 1627 11339
rect 1627 11305 1636 11339
rect 1584 11296 1636 11305
rect 5356 11228 5408 11280
rect 1768 11135 1820 11144
rect 1768 11101 1777 11135
rect 1777 11101 1811 11135
rect 1811 11101 1820 11135
rect 1768 11092 1820 11101
rect 2044 11135 2096 11144
rect 2044 11101 2078 11135
rect 2078 11101 2096 11135
rect 2044 11092 2096 11101
rect 3148 11092 3200 11144
rect 5264 11092 5316 11144
rect 2136 11024 2188 11076
rect 2780 10956 2832 11008
rect 4620 10956 4672 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 2228 10752 2280 10804
rect 1768 10684 1820 10736
rect 2412 10548 2464 10600
rect 3424 10684 3476 10736
rect 5264 10752 5316 10804
rect 2780 10591 2832 10600
rect 2780 10557 2789 10591
rect 2789 10557 2823 10591
rect 2823 10557 2832 10591
rect 2780 10548 2832 10557
rect 3056 10591 3108 10600
rect 3056 10557 3065 10591
rect 3065 10557 3099 10591
rect 3099 10557 3108 10591
rect 3056 10548 3108 10557
rect 2964 10412 3016 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 3056 10208 3108 10260
rect 3148 10072 3200 10124
rect 4712 10115 4764 10124
rect 4712 10081 4721 10115
rect 4721 10081 4755 10115
rect 4755 10081 4764 10115
rect 4712 10072 4764 10081
rect 2780 10004 2832 10056
rect 1400 9936 1452 9988
rect 1768 9936 1820 9988
rect 2504 9979 2556 9988
rect 2504 9945 2513 9979
rect 2513 9945 2547 9979
rect 2547 9945 2556 9979
rect 2504 9936 2556 9945
rect 2964 9936 3016 9988
rect 4620 9936 4672 9988
rect 3332 9911 3384 9920
rect 3332 9877 3341 9911
rect 3341 9877 3375 9911
rect 3375 9877 3384 9911
rect 3332 9868 3384 9877
rect 3424 9911 3476 9920
rect 3424 9877 3433 9911
rect 3433 9877 3467 9911
rect 3467 9877 3476 9911
rect 3424 9868 3476 9877
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 2504 9664 2556 9716
rect 2688 9639 2740 9648
rect 2688 9605 2697 9639
rect 2697 9605 2731 9639
rect 2731 9605 2740 9639
rect 2688 9596 2740 9605
rect 2412 9571 2464 9580
rect 2412 9537 2421 9571
rect 2421 9537 2455 9571
rect 2455 9537 2464 9571
rect 2412 9528 2464 9537
rect 3332 9528 3384 9580
rect 3424 9460 3476 9512
rect 2964 9392 3016 9444
rect 3056 9324 3108 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 3056 9163 3108 9172
rect 3056 9129 3065 9163
rect 3065 9129 3099 9163
rect 3099 9129 3108 9163
rect 3056 9120 3108 9129
rect 3332 9052 3384 9104
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 2964 8916 3016 8968
rect 5264 8916 5316 8968
rect 3240 8891 3292 8900
rect 3240 8857 3249 8891
rect 3249 8857 3283 8891
rect 3283 8857 3292 8891
rect 3240 8848 3292 8857
rect 3424 8891 3476 8900
rect 3424 8857 3433 8891
rect 3433 8857 3467 8891
rect 3467 8857 3476 8891
rect 3424 8848 3476 8857
rect 3608 8891 3660 8900
rect 3608 8857 3617 8891
rect 3617 8857 3651 8891
rect 3651 8857 3660 8891
rect 3608 8848 3660 8857
rect 4620 8780 4672 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 5264 8576 5316 8628
rect 1400 8440 1452 8492
rect 3056 8415 3108 8424
rect 3056 8381 3065 8415
rect 3065 8381 3099 8415
rect 3099 8381 3108 8415
rect 3056 8372 3108 8381
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 3056 8032 3108 8084
rect 4712 7896 4764 7948
rect 3608 7828 3660 7880
rect 4620 7828 4672 7880
rect 5264 7828 5316 7880
rect 5816 7692 5868 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 2964 7284 3016 7336
rect 3240 7216 3292 7268
rect 3516 7191 3568 7200
rect 3516 7157 3525 7191
rect 3525 7157 3559 7191
rect 3559 7157 3568 7191
rect 3516 7148 3568 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 3240 6808 3292 6860
rect 2044 6672 2096 6724
rect 3424 6740 3476 6792
rect 2964 6715 3016 6724
rect 2964 6681 2973 6715
rect 2973 6681 3007 6715
rect 3007 6681 3016 6715
rect 2964 6672 3016 6681
rect 4620 6672 4672 6724
rect 2780 6647 2832 6656
rect 2780 6613 2789 6647
rect 2789 6613 2823 6647
rect 2823 6613 2832 6647
rect 2780 6604 2832 6613
rect 3056 6647 3108 6656
rect 3056 6613 3065 6647
rect 3065 6613 3099 6647
rect 3099 6613 3108 6647
rect 3056 6604 3108 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 2044 6443 2096 6452
rect 2044 6409 2053 6443
rect 2053 6409 2087 6443
rect 2087 6409 2096 6443
rect 2044 6400 2096 6409
rect 1400 6332 1452 6384
rect 2688 6332 2740 6384
rect 3056 6264 3108 6316
rect 3516 6332 3568 6384
rect 2964 6196 3016 6248
rect 2780 6128 2832 6180
rect 4620 6060 4672 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 3608 5695 3660 5704
rect 3608 5661 3617 5695
rect 3617 5661 3651 5695
rect 3651 5661 3660 5695
rect 3608 5652 3660 5661
rect 5356 5652 5408 5704
rect 2964 5559 3016 5568
rect 2964 5525 2973 5559
rect 2973 5525 3007 5559
rect 3007 5525 3016 5559
rect 2964 5516 3016 5525
rect 4712 5516 4764 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 2964 5312 3016 5364
rect 2688 5244 2740 5296
rect 2780 5176 2832 5228
rect 3976 5219 4028 5228
rect 3976 5185 4010 5219
rect 4010 5185 4028 5219
rect 3976 5176 4028 5185
rect 2504 4972 2556 5024
rect 4804 4972 4856 5024
rect 5356 4972 5408 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 3976 4768 4028 4820
rect 4712 4675 4764 4684
rect 4712 4641 4721 4675
rect 4721 4641 4755 4675
rect 4755 4641 4764 4675
rect 4712 4632 4764 4641
rect 4804 4675 4856 4684
rect 4804 4641 4813 4675
rect 4813 4641 4847 4675
rect 4847 4641 4856 4675
rect 4804 4632 4856 4641
rect 4620 4607 4672 4616
rect 4620 4573 4629 4607
rect 4629 4573 4663 4607
rect 4663 4573 4672 4607
rect 4620 4564 4672 4573
rect 2504 4539 2556 4548
rect 2504 4505 2538 4539
rect 2538 4505 2556 4539
rect 2504 4496 2556 4505
rect 2688 4496 2740 4548
rect 3608 4471 3660 4480
rect 3608 4437 3617 4471
rect 3617 4437 3651 4471
rect 3651 4437 3660 4471
rect 3608 4428 3660 4437
rect 4160 4428 4212 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 4160 4088 4212 4140
rect 5264 3952 5316 4004
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 5356 2388 5408 2440
rect 6368 2252 6420 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 5262 22400 5318 22409
rect 5262 22335 5318 22344
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 5276 21690 5304 22335
rect 5264 21684 5316 21690
rect 5264 21626 5316 21632
rect 4804 21548 4856 21554
rect 4804 21490 4856 21496
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4816 21010 4844 21490
rect 4804 21004 4856 21010
rect 4804 20946 4856 20952
rect 4620 20800 4672 20806
rect 4620 20742 4672 20748
rect 2504 20460 2556 20466
rect 2504 20402 2556 20408
rect 3700 20460 3752 20466
rect 3700 20402 3752 20408
rect 3976 20460 4028 20466
rect 3976 20402 4028 20408
rect 2516 20058 2544 20402
rect 3608 20256 3660 20262
rect 3608 20198 3660 20204
rect 2504 20052 2556 20058
rect 2504 19994 2556 20000
rect 3620 19922 3648 20198
rect 3608 19916 3660 19922
rect 3608 19858 3660 19864
rect 2780 19848 2832 19854
rect 2780 19790 2832 19796
rect 2872 19848 2924 19854
rect 2872 19790 2924 19796
rect 2792 19378 2820 19790
rect 2884 19514 2912 19790
rect 2964 19712 3016 19718
rect 2964 19654 3016 19660
rect 2976 19514 3004 19654
rect 2872 19508 2924 19514
rect 2872 19450 2924 19456
rect 2964 19508 3016 19514
rect 2964 19450 3016 19456
rect 2780 19372 2832 19378
rect 2780 19314 2832 19320
rect 3148 19372 3200 19378
rect 3148 19314 3200 19320
rect 2320 19304 2372 19310
rect 2320 19246 2372 19252
rect 2332 18970 2360 19246
rect 2320 18964 2372 18970
rect 2320 18906 2372 18912
rect 1676 18760 1728 18766
rect 1676 18702 1728 18708
rect 1688 18290 1716 18702
rect 1676 18284 1728 18290
rect 1676 18226 1728 18232
rect 1688 17814 1716 18226
rect 1676 17808 1728 17814
rect 662 17776 718 17785
rect 1676 17750 1728 17756
rect 662 17711 718 17720
rect 676 17678 704 17711
rect 664 17672 716 17678
rect 664 17614 716 17620
rect 2228 16788 2280 16794
rect 2228 16730 2280 16736
rect 2136 16652 2188 16658
rect 2136 16594 2188 16600
rect 1952 16108 2004 16114
rect 1952 16050 2004 16056
rect 1964 15162 1992 16050
rect 2044 15904 2096 15910
rect 2044 15846 2096 15852
rect 2056 15434 2084 15846
rect 2044 15428 2096 15434
rect 2044 15370 2096 15376
rect 1952 15156 2004 15162
rect 1952 15098 2004 15104
rect 2148 15042 2176 16594
rect 2240 16114 2268 16730
rect 2332 16658 2360 18906
rect 2780 18760 2832 18766
rect 2780 18702 2832 18708
rect 2792 18426 2820 18702
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 2792 17678 2820 18362
rect 3056 18352 3108 18358
rect 3056 18294 3108 18300
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 3068 17202 3096 18294
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 2320 16652 2372 16658
rect 2320 16594 2372 16600
rect 2228 16108 2280 16114
rect 2228 16050 2280 16056
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 2056 15026 2176 15042
rect 2044 15020 2176 15026
rect 2096 15014 2176 15020
rect 2044 14962 2096 14968
rect 2056 11898 2084 14962
rect 2516 14618 2544 16050
rect 3068 15502 3096 17138
rect 3160 16590 3188 19314
rect 3712 18290 3740 20402
rect 3988 19514 4016 20402
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4632 19786 4660 20742
rect 4816 20602 4844 20946
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4804 20596 4856 20602
rect 4804 20538 4856 20544
rect 5264 19916 5316 19922
rect 5264 19858 5316 19864
rect 4620 19780 4672 19786
rect 4620 19722 4672 19728
rect 4344 19712 4396 19718
rect 4344 19654 4396 19660
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 4356 19310 4384 19654
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 4988 19508 5040 19514
rect 4988 19450 5040 19456
rect 5000 19417 5028 19450
rect 4986 19408 5042 19417
rect 4804 19372 4856 19378
rect 4986 19343 5042 19352
rect 4804 19314 4856 19320
rect 4344 19304 4396 19310
rect 4344 19246 4396 19252
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4068 18624 4120 18630
rect 4068 18566 4120 18572
rect 4080 18358 4108 18566
rect 4068 18352 4120 18358
rect 4068 18294 4120 18300
rect 3700 18284 3752 18290
rect 3700 18226 3752 18232
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17746 4660 18022
rect 4724 17882 4752 18702
rect 4816 18426 4844 19314
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 4712 17876 4764 17882
rect 4712 17818 4764 17824
rect 5276 17746 5304 19858
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 4712 17740 4764 17746
rect 4712 17682 4764 17688
rect 5264 17740 5316 17746
rect 5264 17682 5316 17688
rect 4068 17536 4120 17542
rect 4068 17478 4120 17484
rect 3332 17196 3384 17202
rect 3332 17138 3384 17144
rect 3344 16794 3372 17138
rect 4080 16998 4108 17478
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 4080 16658 4108 16934
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 3884 16652 3936 16658
rect 3884 16594 3936 16600
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 3148 16584 3200 16590
rect 3148 16526 3200 16532
rect 3160 15706 3188 16526
rect 3148 15700 3200 15706
rect 3148 15642 3200 15648
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 3700 15496 3752 15502
rect 3700 15438 3752 15444
rect 2596 15428 2648 15434
rect 2596 15370 2648 15376
rect 3516 15428 3568 15434
rect 3516 15370 3568 15376
rect 2608 15026 2636 15370
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 3332 15360 3384 15366
rect 3332 15302 3384 15308
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 2688 15020 2740 15026
rect 2688 14962 2740 14968
rect 2504 14612 2556 14618
rect 2504 14554 2556 14560
rect 2608 14346 2636 14962
rect 2136 14340 2188 14346
rect 2136 14282 2188 14288
rect 2596 14340 2648 14346
rect 2596 14282 2648 14288
rect 2148 12850 2176 14282
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2240 12986 2268 13126
rect 2228 12980 2280 12986
rect 2228 12922 2280 12928
rect 2136 12844 2188 12850
rect 2136 12786 2188 12792
rect 2596 12844 2648 12850
rect 2596 12786 2648 12792
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 1584 11824 1636 11830
rect 1584 11766 1636 11772
rect 1596 11354 1624 11766
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 2056 11150 2084 11494
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 2044 11144 2096 11150
rect 2044 11086 2096 11092
rect 1780 10742 1808 11086
rect 2148 11082 2176 12786
rect 2412 12640 2464 12646
rect 2412 12582 2464 12588
rect 2424 12170 2452 12582
rect 2412 12164 2464 12170
rect 2412 12106 2464 12112
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 2136 11076 2188 11082
rect 2136 11018 2188 11024
rect 2240 10810 2268 11494
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 1768 10736 1820 10742
rect 1768 10678 1820 10684
rect 1780 9994 1808 10678
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 1400 9988 1452 9994
rect 1400 9930 1452 9936
rect 1768 9988 1820 9994
rect 1768 9930 1820 9936
rect 1412 8974 1440 9930
rect 2424 9586 2452 10542
rect 2504 9988 2556 9994
rect 2504 9930 2556 9936
rect 2516 9722 2544 9930
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1412 8498 1440 8910
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 6866 1440 8434
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1412 6390 1440 6802
rect 2044 6724 2096 6730
rect 2044 6666 2096 6672
rect 2056 6458 2084 6666
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 1400 6384 1452 6390
rect 1400 6326 1452 6332
rect 2608 5817 2636 12786
rect 2700 12646 2728 14962
rect 2792 14958 2820 15302
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2792 14550 2820 14894
rect 2780 14544 2832 14550
rect 2780 14486 2832 14492
rect 2884 14346 2912 15098
rect 3344 14550 3372 15302
rect 3528 15162 3556 15370
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 3712 14822 3740 15438
rect 3896 15366 3924 16594
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 3884 15360 3936 15366
rect 3884 15302 3936 15308
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3332 14544 3384 14550
rect 3332 14486 3384 14492
rect 2872 14340 2924 14346
rect 2872 14282 2924 14288
rect 2884 13394 2912 14282
rect 3712 13870 3740 14758
rect 3988 14618 4016 15438
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 4080 14006 4108 15302
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4724 14482 4752 17682
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4068 14000 4120 14006
rect 4068 13942 4120 13948
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 3700 13864 3752 13870
rect 3700 13806 3752 13812
rect 2872 13388 2924 13394
rect 2872 13330 2924 13336
rect 2884 13002 2912 13330
rect 2884 12974 3004 13002
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2700 9654 2728 12582
rect 2884 12442 2912 12854
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 2872 12300 2924 12306
rect 2872 12242 2924 12248
rect 2884 11898 2912 12242
rect 2976 12102 3004 12974
rect 3068 12238 3096 13806
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4620 13456 4672 13462
rect 4620 13398 4672 13404
rect 4436 13184 4488 13190
rect 4436 13126 4488 13132
rect 4448 12986 4476 13126
rect 4436 12980 4488 12986
rect 4436 12922 4488 12928
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 12306 4660 13398
rect 4724 13394 4752 14418
rect 4816 14278 4844 16526
rect 5264 16448 5316 16454
rect 5262 16416 5264 16425
rect 5316 16416 5318 16425
rect 4874 16348 5182 16357
rect 5262 16351 5318 16360
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 4816 14074 4844 14214
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4896 13456 4948 13462
rect 4894 13424 4896 13433
rect 4948 13424 4950 13433
rect 4712 13388 4764 13394
rect 4894 13359 4950 13368
rect 4712 13330 4764 13336
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 3068 11762 3096 12174
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 3160 11150 3188 12174
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 2792 10606 2820 10950
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 2792 10062 2820 10542
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2976 9994 3004 10406
rect 3068 10266 3096 10542
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 3160 10130 3188 11086
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 2688 9648 2740 9654
rect 2688 9590 2740 9596
rect 2976 9450 3004 9930
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2976 8974 3004 9386
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 3068 9178 3096 9318
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2976 7342 3004 8910
rect 3252 8906 3280 11834
rect 3896 11830 3924 12038
rect 3884 11824 3936 11830
rect 3884 11766 3936 11772
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4620 11008 4672 11014
rect 4620 10950 4672 10956
rect 3424 10736 3476 10742
rect 3424 10678 3476 10684
rect 3436 9926 3464 10678
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4632 9994 4660 10950
rect 4724 10130 4752 13330
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4816 12782 4844 13262
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4816 11898 4844 12718
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 5356 11280 5408 11286
rect 5356 11222 5408 11228
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 5276 10810 5304 11086
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5368 10441 5396 11222
rect 5354 10432 5410 10441
rect 5354 10367 5410 10376
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 3332 9920 3384 9926
rect 3332 9862 3384 9868
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3344 9586 3372 9862
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3344 9110 3372 9522
rect 3436 9518 3464 9862
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3436 8906 3464 9454
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 3240 8900 3292 8906
rect 3240 8842 3292 8848
rect 3424 8900 3476 8906
rect 3424 8842 3476 8848
rect 3608 8900 3660 8906
rect 3608 8842 3660 8848
rect 3056 8424 3108 8430
rect 3056 8366 3108 8372
rect 3068 8090 3096 8366
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 2976 6730 3004 7278
rect 3252 7274 3280 8842
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3252 6866 3280 7210
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 3436 6798 3464 8842
rect 3620 7886 3648 8842
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7886 4660 8774
rect 4724 7954 4752 10066
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5276 8634 5304 8910
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2688 6384 2740 6390
rect 2688 6326 2740 6332
rect 2594 5808 2650 5817
rect 2594 5743 2650 5752
rect 2700 5302 2728 6326
rect 2792 6186 2820 6598
rect 2976 6254 3004 6666
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 3068 6322 3096 6598
rect 3528 6390 3556 7142
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4724 6914 4752 7890
rect 5276 7886 5304 8570
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 5828 7449 5856 7686
rect 5814 7440 5870 7449
rect 5814 7375 5870 7384
rect 4724 6886 4844 6914
rect 4620 6724 4672 6730
rect 4620 6666 4672 6672
rect 3516 6384 3568 6390
rect 3516 6326 3568 6332
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 2780 6180 2832 6186
rect 2780 6122 2832 6128
rect 2688 5296 2740 5302
rect 2688 5238 2740 5244
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 2516 4554 2544 4966
rect 2700 4554 2728 5238
rect 2792 5234 2820 6122
rect 4632 6118 4660 6666
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 3608 5704 3660 5710
rect 3608 5646 3660 5652
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2976 5370 3004 5510
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 2504 4548 2556 4554
rect 2504 4490 2556 4496
rect 2688 4548 2740 4554
rect 2688 4490 2740 4496
rect 3620 4486 3648 5646
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 3988 4826 4016 5170
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 4632 4622 4660 6054
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4724 4690 4752 5510
rect 4816 5030 4844 6886
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5368 5030 5396 5646
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 4816 4690 4844 4966
rect 4712 4684 4764 4690
rect 4712 4626 4764 4632
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 3608 4480 3660 4486
rect 3608 4422 3660 4428
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 5262 4448 5318 4457
rect 4172 4146 4200 4422
rect 4874 4380 5182 4389
rect 5262 4383 5318 4392
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 5276 4010 5304 4383
rect 5264 4004 5316 4010
rect 5264 3946 5316 3952
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 5368 2446 5396 4966
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 6368 2304 6420 2310
rect 6368 2246 6420 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 6380 1465 6408 2246
rect 6366 1456 6422 1465
rect 6366 1391 6422 1400
<< via2 >>
rect 5262 22344 5318 22400
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 662 17720 718 17776
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4986 19352 5042 19408
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 5262 16396 5264 16416
rect 5264 16396 5316 16416
rect 5316 16396 5318 16416
rect 5262 16360 5318 16396
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4894 13404 4896 13424
rect 4896 13404 4948 13424
rect 4948 13404 4950 13424
rect 4894 13368 4950 13404
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 5354 10376 5410 10432
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 2594 5752 2650 5808
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 5814 7384 5870 7440
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 5262 4392 5318 4448
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 6366 1400 6422 1456
<< metal3 >>
rect 5257 22402 5323 22405
rect 6540 22402 6600 22432
rect 5257 22400 6600 22402
rect 5257 22344 5262 22400
rect 5318 22344 6600 22400
rect 5257 22342 6600 22344
rect 5257 22339 5323 22342
rect 6540 22312 6600 22342
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 4981 19410 5047 19413
rect 6540 19410 6600 19440
rect 4981 19408 6600 19410
rect 4981 19352 4986 19408
rect 5042 19352 6600 19408
rect 4981 19350 6600 19352
rect 4981 19347 5047 19350
rect 6540 19320 6600 19350
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 0 17778 60 17808
rect 657 17778 723 17781
rect 0 17776 723 17778
rect 0 17720 662 17776
rect 718 17720 723 17776
rect 0 17718 723 17720
rect 0 17688 60 17718
rect 657 17715 723 17718
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 5257 16418 5323 16421
rect 6540 16418 6600 16448
rect 5257 16416 6600 16418
rect 5257 16360 5262 16416
rect 5318 16360 6600 16416
rect 5257 16358 6600 16360
rect 5257 16355 5323 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 6540 16328 6600 16358
rect 4870 16287 5186 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 4889 13426 4955 13429
rect 6540 13426 6600 13456
rect 4889 13424 6600 13426
rect 4889 13368 4894 13424
rect 4950 13368 6600 13424
rect 4889 13366 6600 13368
rect 4889 13363 4955 13366
rect 6540 13336 6600 13366
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 5349 10434 5415 10437
rect 6540 10434 6600 10464
rect 5349 10432 6600 10434
rect 5349 10376 5354 10432
rect 5410 10376 6600 10432
rect 5349 10374 6600 10376
rect 5349 10371 5415 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 6540 10344 6600 10374
rect 4210 10303 4526 10304
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 5809 7442 5875 7445
rect 6540 7442 6600 7472
rect 5809 7440 6600 7442
rect 5809 7384 5814 7440
rect 5870 7384 6600 7440
rect 5809 7382 6600 7384
rect 5809 7379 5875 7382
rect 6540 7352 6600 7382
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 0 5810 60 5840
rect 2589 5810 2655 5813
rect 0 5808 2655 5810
rect 0 5752 2594 5808
rect 2650 5752 2655 5808
rect 0 5750 2655 5752
rect 0 5720 60 5750
rect 2589 5747 2655 5750
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 5257 4450 5323 4453
rect 6540 4450 6600 4480
rect 5257 4448 6600 4450
rect 5257 4392 5262 4448
rect 5318 4392 6600 4448
rect 5257 4390 6600 4392
rect 5257 4387 5323 4390
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 6540 4360 6600 4390
rect 4870 4319 5186 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 6361 1458 6427 1461
rect 6540 1458 6600 1488
rect 6361 1456 6600 1458
rect 6361 1400 6366 1456
rect 6422 1400 6600 1456
rect 6361 1398 6600 1400
rect 6361 1395 6427 1398
rect 6540 1368 6600 1398
<< via3 >>
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 21248 4528 21808
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 21792 5188 21808
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__nand2b_2  _31_
timestamp -3599
transform 1 0 1840 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _32_
timestamp -3599
transform 1 0 3036 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _33_
timestamp -3599
transform -1 0 3404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _34_
timestamp -3599
transform 1 0 2024 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _35_
timestamp -3599
transform -1 0 2668 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _36_
timestamp -3599
transform -1 0 3680 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _37_
timestamp -3599
transform -1 0 3312 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _38_
timestamp -3599
transform 1 0 2300 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _39_
timestamp -3599
transform -1 0 3680 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _40_
timestamp 1562532584
transform -1 0 1748 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _41_
timestamp -3599
transform -1 0 2484 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _42_
timestamp -3599
transform -1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _43_
timestamp -3599
transform -1 0 2484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _44_
timestamp -3599
transform 1 0 2116 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _45_
timestamp -3599
transform -1 0 2944 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _46_
timestamp -3599
transform 1 0 1840 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _47_
timestamp -3599
transform 1 0 2024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _48_
timestamp -3599
transform -1 0 3588 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _49_
timestamp -3599
transform -1 0 3128 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _50_
timestamp -3599
transform -1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _51_
timestamp -3599
transform -1 0 3312 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _52_
timestamp -3599
transform 1 0 2392 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_4  _53_
timestamp -3599
transform -1 0 3220 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_1  _54_
timestamp -3599
transform 1 0 4232 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _55_
timestamp -3599
transform 1 0 2760 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _56_
timestamp -3599
transform 1 0 3956 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _57_
timestamp -3599
transform 1 0 4048 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _58_
timestamp -3599
transform 1 0 3772 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _59_
timestamp -3599
transform 1 0 4048 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _60_
timestamp -3599
transform 1 0 4140 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _61_
timestamp -3599
transform 1 0 4048 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _62_
timestamp -3599
transform 1 0 3404 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _63_
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _64_
timestamp -3599
transform 1 0 1380 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _65_
timestamp -3599
transform 1 0 1748 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _66_
timestamp -3599
transform 1 0 1472 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _67_
timestamp -3599
transform 1 0 1380 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _68_
timestamp -3599
transform 1 0 3036 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _69_
timestamp -3599
transform 1 0 2208 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _70_
timestamp -3599
transform 1 0 3680 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _71_
timestamp -3599
transform 1 0 2208 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _72_
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _73_
timestamp -3599
transform 1 0 3680 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _74_
timestamp -3599
transform 1 0 3588 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _75_
timestamp -3599
transform 1 0 3680 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _76_
timestamp -3599
transform 1 0 3680 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _77_
timestamp -3599
transform 1 0 3680 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _78_
timestamp -3599
transform 1 0 1380 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp -3599
transform 1 0 2576 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp -3599
transform 1 0 2668 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp -3599
transform 1 0 2668 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  clkload0
timestamp -3599
transform 1 0 2392 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3
timestamp -3599
transform 1 0 1380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11
timestamp -3599
transform 1 0 2116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19
timestamp -3599
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29
timestamp -3599
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37
timestamp -3599
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3
timestamp -3599
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_11
timestamp -3599
transform 1 0 2116 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_19
timestamp -3599
transform 1 0 2852 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_27
timestamp -3599
transform 1 0 3588 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_35
timestamp -3599
transform 1 0 4324 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_43
timestamp -3599
transform 1 0 5060 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp -3599
transform 1 0 1380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_11
timestamp -3599
transform 1 0 2116 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_19
timestamp -3599
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_29
timestamp -3599
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_37
timestamp -3599
transform 1 0 4508 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_43
timestamp -3599
transform 1 0 5060 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp -3599
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_11
timestamp -3599
transform 1 0 2116 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_19
timestamp -3599
transform 1 0 2852 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_27
timestamp -3599
transform 1 0 3588 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_35
timestamp -3599
transform 1 0 4324 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_39
timestamp -3599
transform 1 0 4692 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp -3599
transform 1 0 1380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_11
timestamp -3599
transform 1 0 2116 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp -3599
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_33
timestamp -3599
transform 1 0 4140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_43
timestamp -3599
transform 1 0 5060 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3
timestamp -3599
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_11
timestamp -3599
transform 1 0 2116 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_17
timestamp -3599
transform 1 0 2668 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_27
timestamp -3599
transform 1 0 3588 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp -3599
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_11
timestamp -3599
transform 1 0 2116 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_19
timestamp -3599
transform 1 0 2852 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_29
timestamp -3599
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_35
timestamp -3599
transform 1 0 4324 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp -3599
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_9
timestamp -3599
transform 1 0 1932 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_16
timestamp -3599
transform 1 0 2576 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_24
timestamp -3599
transform 1 0 3312 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_41
timestamp -3599
transform 1 0 4876 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp -3599
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_29
timestamp -3599
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_37
timestamp -3599
transform 1 0 4508 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_43
timestamp -3599
transform 1 0 5060 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp -3599
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_11
timestamp -3599
transform 1 0 2116 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_19
timestamp -3599
transform 1 0 2852 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_27
timestamp -3599
transform 1 0 3588 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_35
timestamp -3599
transform 1 0 4324 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_43
timestamp -3599
transform 1 0 5060 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_11
timestamp -3599
transform 1 0 2116 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp -3599
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp -3599
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp -3599
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_11
timestamp -3599
transform 1 0 2116 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_19
timestamp -3599
transform 1 0 2852 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_29
timestamp -3599
transform 1 0 3772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_35
timestamp -3599
transform 1 0 4324 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3
timestamp -3599
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_37
timestamp -3599
transform 1 0 4508 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_43
timestamp -3599
transform 1 0 5060 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp -3599
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_11
timestamp -3599
transform 1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_29
timestamp -3599
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_41
timestamp -3599
transform 1 0 4876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_3
timestamp -3599
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_11
timestamp -3599
transform 1 0 2116 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp -3599
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp -3599
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp -3599
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_29
timestamp -3599
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp -3599
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp -3599
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_15
timestamp -3599
transform 1 0 2484 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_23
timestamp -3599
transform 1 0 3220 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_43
timestamp -3599
transform 1 0 5060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp -3599
transform 1 0 1380 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp -3599
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_29
timestamp -3599
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_38
timestamp -3599
transform 1 0 4600 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp -3599
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_15
timestamp -3599
transform 1 0 2484 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp -3599
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_11
timestamp -3599
transform 1 0 2116 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_15
timestamp -3599
transform 1 0 2484 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp -3599
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_38
timestamp -3599
transform 1 0 4600 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp -3599
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_11
timestamp -3599
transform 1 0 2116 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_19
timestamp -3599
transform 1 0 2852 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_27
timestamp -3599
transform 1 0 3588 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp -3599
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_11
timestamp -3599
transform 1 0 2116 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_29
timestamp -3599
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_41
timestamp -3599
transform 1 0 4876 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp -3599
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp -3599
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_37
timestamp -3599
transform 1 0 4508 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_43
timestamp -3599
transform 1 0 5060 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_19
timestamp -3599
transform 1 0 2852 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp -3599
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_29
timestamp -3599
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_40
timestamp -3599
transform 1 0 4784 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp -3599
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_9
timestamp -3599
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_13
timestamp -3599
transform 1 0 2300 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_21
timestamp -3599
transform 1 0 3036 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_29
timestamp -3599
transform 1 0 3772 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_37
timestamp -3599
transform 1 0 4508 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_43
timestamp -3599
transform 1 0 5060 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp -3599
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_11
timestamp -3599
transform 1 0 2116 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_17
timestamp -3599
transform 1 0 2668 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_25
timestamp -3599
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_37
timestamp -3599
transform 1 0 4508 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp -3599
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_11
timestamp -3599
transform 1 0 2116 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_19
timestamp -3599
transform 1 0 2852 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_37
timestamp -3599
transform 1 0 4508 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_43
timestamp -3599
transform 1 0 5060 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_6
timestamp -3599
transform 1 0 1656 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_23
timestamp -3599
transform 1 0 3220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp -3599
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_29
timestamp -3599
transform 1 0 3772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_42
timestamp -3599
transform 1 0 4968 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_19
timestamp -3599
transform 1 0 2852 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp -3599
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_7
timestamp -3599
transform 1 0 1748 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_15
timestamp -3599
transform 1 0 2484 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_23
timestamp -3599
transform 1 0 3220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp -3599
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_29
timestamp -3599
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_40
timestamp -3599
transform 1 0 4784 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_3
timestamp -3599
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_11
timestamp -3599
transform 1 0 2116 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_17
timestamp -3599
transform 1 0 2668 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_24
timestamp -3599
transform 1 0 3312 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_3
timestamp -3599
transform 1 0 1380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_11
timestamp -3599
transform 1 0 2116 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_29
timestamp -3599
transform 1 0 3772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_41
timestamp -3599
transform 1 0 4876 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_3
timestamp -3599
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_11
timestamp -3599
transform 1 0 2116 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_3
timestamp -3599
transform 1 0 1380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_11
timestamp -3599
transform 1 0 2116 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_19
timestamp -3599
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp -3599
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_29
timestamp -3599
transform 1 0 3772 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_35
timestamp -3599
transform 1 0 4324 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_3
timestamp -3599
transform 1 0 1380 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_11
timestamp -3599
transform 1 0 2116 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_19
timestamp -3599
transform 1 0 2852 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_27
timestamp -3599
transform 1 0 3588 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_29
timestamp -3599
transform 1 0 3772 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_37
timestamp -3599
transform 1 0 4508 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp -3599
transform -1 0 5152 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp -3599
transform 1 0 2944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp -3599
transform -1 0 5152 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp -3599
transform 1 0 2944 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp -3599
transform 1 0 2944 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp -3599
transform -1 0 4784 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp -3599
transform -1 0 5152 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp -3599
transform -1 0 4784 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp -3599
transform -1 0 3680 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp -3599
transform -1 0 5152 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp -3599
transform -1 0 4600 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp -3599
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp -3599
transform -1 0 4784 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp -3599
transform -1 0 5152 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp -3599
transform -1 0 3680 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp -3599
transform -1 0 4508 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp -3599
transform -1 0 3312 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp -3599
transform 1 0 1380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output2
timestamp -3599
transform -1 0 5152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp -3599
transform 1 0 4784 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp -3599
transform 1 0 4784 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp -3599
transform -1 0 4416 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp -3599
transform -1 0 5152 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp -3599
transform 1 0 4784 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp -3599
transform 1 0 4784 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp -3599
transform 1 0 4784 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_36
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 5428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_37
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 5428 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_38
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 5428 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_39
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 5428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_40
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 5428 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_41
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 5428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_42
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 5428 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_43
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 5428 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_44
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 5428 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_45
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 5428 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_46
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 5428 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_47
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 5428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_48
timestamp -3599
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -3599
transform -1 0 5428 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_49
timestamp -3599
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -3599
transform -1 0 5428 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_50
timestamp -3599
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -3599
transform -1 0 5428 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_51
timestamp -3599
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -3599
transform -1 0 5428 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_52
timestamp -3599
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -3599
transform -1 0 5428 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_53
timestamp -3599
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -3599
transform -1 0 5428 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_54
timestamp -3599
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp -3599
transform -1 0 5428 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_55
timestamp -3599
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp -3599
transform -1 0 5428 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_56
timestamp -3599
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp -3599
transform -1 0 5428 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_57
timestamp -3599
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp -3599
transform -1 0 5428 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_58
timestamp -3599
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp -3599
transform -1 0 5428 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_59
timestamp -3599
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp -3599
transform -1 0 5428 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_60
timestamp -3599
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp -3599
transform -1 0 5428 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_61
timestamp -3599
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp -3599
transform -1 0 5428 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_62
timestamp -3599
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp -3599
transform -1 0 5428 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_63
timestamp -3599
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp -3599
transform -1 0 5428 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_64
timestamp -3599
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp -3599
transform -1 0 5428 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_65
timestamp -3599
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp -3599
transform -1 0 5428 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_66
timestamp -3599
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp -3599
transform -1 0 5428 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_67
timestamp -3599
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp -3599
transform -1 0 5428 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_68
timestamp -3599
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp -3599
transform -1 0 5428 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_69
timestamp -3599
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp -3599
transform -1 0 5428 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_70
timestamp -3599
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp -3599
transform -1 0 5428 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_71
timestamp -3599
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp -3599
transform -1 0 5428 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_73
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_74
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_75
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_76
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_77
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_78
timestamp -3599
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_79
timestamp -3599
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_80
timestamp -3599
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_81
timestamp -3599
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_82
timestamp -3599
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_83
timestamp -3599
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_84
timestamp -3599
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_85
timestamp -3599
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_86
timestamp -3599
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_87
timestamp -3599
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_88
timestamp -3599
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_89
timestamp -3599
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_90
timestamp -3599
transform 1 0 3680 0 -1 21760
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 5720 60 5840 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 6540 1368 6600 1488 0 FreeSans 480 0 0 0 counter_out[0]
port 3 nsew signal output
flabel metal3 s 6540 4360 6600 4480 0 FreeSans 480 0 0 0 counter_out[1]
port 4 nsew signal output
flabel metal3 s 6540 7352 6600 7472 0 FreeSans 480 0 0 0 counter_out[2]
port 5 nsew signal output
flabel metal3 s 6540 10344 6600 10464 0 FreeSans 480 0 0 0 counter_out[3]
port 6 nsew signal output
flabel metal3 s 6540 13336 6600 13456 0 FreeSans 480 0 0 0 counter_out[4]
port 7 nsew signal output
flabel metal3 s 6540 16328 6600 16448 0 FreeSans 480 0 0 0 counter_out[5]
port 8 nsew signal output
flabel metal3 s 6540 19320 6600 19440 0 FreeSans 480 0 0 0 counter_out[6]
port 9 nsew signal output
flabel metal3 s 6540 22312 6600 22432 0 FreeSans 480 0 0 0 counter_out[7]
port 10 nsew signal output
flabel metal3 s 0 17688 60 17808 0 FreeSans 480 0 0 0 trigger
port 11 nsew signal input
rlabel metal1 3266 21760 3266 21760 0 VGND
rlabel metal1 3266 21216 3266 21216 0 VPWR
rlabel metal1 3618 6358 3618 6358 0 _00_
rlabel metal2 2070 6562 2070 6562 0 _01_
rlabel metal1 2295 8874 2295 8874 0 _02_
rlabel via1 2065 11118 2065 11118 0 _03_
rlabel metal1 2111 12138 2111 12138 0 _04_
rlabel metal1 1881 15402 1881 15402 0 _05_
rlabel metal2 3358 16966 3358 16966 0 _06_
rlabel metal1 2484 20026 2484 20026 0 _07_
rlabel metal1 4140 4794 4140 4794 0 _08_
rlabel via1 2525 4522 2525 4522 0 _09_
rlabel metal1 3542 8058 3542 8058 0 _10_
rlabel metal1 3588 10234 3588 10234 0 _11_
rlabel metal1 4600 12274 4600 12274 0 _12_
rlabel metal1 4048 14586 4048 14586 0 _13_
rlabel metal1 4462 17850 4462 17850 0 _14_
rlabel metal1 4508 19278 4508 19278 0 _15_
rlabel metal1 3312 6834 3312 6834 0 _16_
rlabel metal1 2668 6290 2668 6290 0 _17_
rlabel metal2 3082 9248 3082 9248 0 _18_
rlabel metal1 3212 8806 3212 8806 0 _19_
rlabel metal1 2300 10778 2300 10778 0 _20_
rlabel metal2 3174 11152 3174 11152 0 _21_
rlabel metal2 1610 11560 1610 11560 0 _22_
rlabel metal1 2990 12410 2990 12410 0 _23_
rlabel metal1 1886 15028 1886 15028 0 _24_
rlabel metal1 2622 16762 2622 16762 0 _25_
rlabel metal2 1978 15606 1978 15606 0 _26_
rlabel metal1 2990 19346 2990 19346 0 _27_
rlabel metal1 3128 16694 3128 16694 0 _28_
rlabel metal2 2990 19584 2990 19584 0 _29_
rlabel metal1 3450 5066 3450 5066 0 _30_
rlabel metal3 1341 5780 1341 5780 0 clk
rlabel metal1 3312 12614 3312 12614 0 clknet_0_clk
rlabel metal1 3450 6324 3450 6324 0 clknet_1_0__leaf_clk
rlabel metal1 2254 20468 2254 20468 0 clknet_1_1__leaf_clk
rlabel metal1 4738 6086 4738 6086 0 counter\[0\]
rlabel metal1 3174 6766 3174 6766 0 counter\[1\]
rlabel metal2 3634 8364 3634 8364 0 counter\[2\]
rlabel metal1 3864 10030 3864 10030 0 counter\[3\]
rlabel metal1 3036 15130 3036 15130 0 counter\[4\]
rlabel metal1 2714 14552 2714 14552 0 counter\[5\]
rlabel metal1 4140 16626 4140 16626 0 counter\[6\]
rlabel metal2 3634 20060 3634 20060 0 counter\[7\]
rlabel metal3 6467 1428 6467 1428 0 counter_out[0]
rlabel metal1 5152 3978 5152 3978 0 counter_out[1]
rlabel metal3 6191 7412 6191 7412 0 counter_out[2]
rlabel metal3 5961 10404 5961 10404 0 counter_out[3]
rlabel metal3 5731 13396 5731 13396 0 counter_out[4]
rlabel metal1 5152 16422 5152 16422 0 counter_out[5]
rlabel metal3 5777 19380 5777 19380 0 counter_out[6]
rlabel metal1 5152 21658 5152 21658 0 counter_out[7]
rlabel metal1 1932 17782 1932 17782 0 net1
rlabel metal1 4554 7854 4554 7854 0 net10
rlabel metal1 3802 8534 3802 8534 0 net11
rlabel metal1 4600 9962 4600 9962 0 net12
rlabel metal1 3802 10710 3802 10710 0 net13
rlabel metal2 4646 17884 4646 17884 0 net14
rlabel metal1 4043 18326 4043 18326 0 net15
rlabel metal1 4600 19754 4600 19754 0 net16
rlabel metal1 4048 19482 4048 19482 0 net17
rlabel metal1 3128 5338 3128 5338 0 net18
rlabel metal2 4462 13056 4462 13056 0 net19
rlabel metal1 5244 4998 5244 4998 0 net2
rlabel via1 3905 11798 3905 11798 0 net20
rlabel metal1 4094 14314 4094 14314 0 net21
rlabel metal1 4043 13974 4043 13974 0 net22
rlabel metal2 4738 5100 4738 5100 0 net23
rlabel metal1 2944 19822 2944 19822 0 net24
rlabel metal1 3450 16490 3450 16490 0 net25
rlabel metal2 2254 13056 2254 13056 0 net26
rlabel metal1 3910 4454 3910 4454 0 net3
rlabel metal1 5198 8602 5198 8602 0 net4
rlabel metal1 5198 11118 5198 11118 0 net5
rlabel metal1 4922 12750 4922 12750 0 net6
rlabel metal1 4968 14042 4968 14042 0 net7
rlabel metal1 4462 18394 4462 18394 0 net8
rlabel metal1 4922 20978 4922 20978 0 net9
rlabel metal3 375 17748 375 17748 0 trigger
rlabel metal2 2806 18564 2806 18564 0 trigger_prev
<< properties >>
string FIXED_BBOX 0 0 6600 24000
<< end >>
