magic
tech sky130A
magscale 1 2
timestamp 1744554176
<< locali >>
rect -4982 11670 -4214 11688
rect -4982 11114 -4950 11670
rect -4394 11114 -4214 11670
rect -4982 10408 -4214 11114
rect 16292 11670 16860 11676
rect 16292 11114 16298 11670
rect 16854 11114 16860 11670
rect 16292 10084 16860 11114
rect 16292 10024 16856 10084
rect 10096 5152 10288 5293
rect 10096 5120 10464 5152
rect 9856 4928 10496 5120
rect 9856 4480 9984 4928
rect 10432 4480 10496 4928
rect 9856 4416 10496 4480
rect 15616 4416 17408 4544
rect 14840 4144 14900 4258
rect 15616 4160 15680 4416
rect 17344 4096 17408 4416
rect 18082 4170 18142 4386
rect 14840 4066 14900 4084
rect 14840 4064 14848 4066
rect 17439 3867 17633 3873
rect 17439 3812 17508 3867
rect 17563 3812 17633 3867
rect 17439 3743 17633 3812
rect -8221 -6953 -7651 -5155
rect -8221 -7511 -8215 -6953
rect -7657 -7511 -7651 -6953
rect -8221 -7517 -7651 -7511
<< viali >>
rect -4950 11114 -4394 11670
rect 16298 11114 16854 11670
rect 9984 4480 10432 4928
rect 14840 4258 14900 4318
rect 18082 4386 18142 4446
rect 17508 3812 17563 3867
rect 15010 3746 15069 3805
rect -8215 -7511 -7657 -6953
<< metal1 >>
rect -4962 11748 -4956 12316
rect -4388 11748 -4382 12316
rect 16286 11748 16292 12316
rect 16860 11748 16866 12316
rect -4956 11670 -4388 11748
rect -4956 11114 -4950 11670
rect -4394 11114 -4388 11670
rect -4956 11102 -4388 11114
rect 16292 11670 16860 11748
rect 16292 11114 16298 11670
rect 16854 11114 16860 11670
rect 16292 11102 16860 11114
rect -14100 4892 -1456 5084
rect 988 3636 2854 3700
rect 3732 3232 3924 5744
rect 9972 4928 10444 4934
rect 9972 4480 9984 4928
rect 10432 4480 10444 4928
rect 19264 4800 19392 6720
rect 9972 4474 10444 4480
rect 14807 4673 19392 4800
rect 9984 4448 10432 4474
rect 14807 4318 14934 4673
rect 14976 4672 19392 4673
rect 18076 4452 18148 4458
rect 18070 4392 18076 4452
rect 18148 4392 18154 4452
rect 18070 4386 18082 4392
rect 18142 4386 18154 4392
rect 18070 4380 18154 4386
rect 14807 4289 14840 4318
rect 14828 4258 14840 4289
rect 14900 4289 14934 4318
rect 14900 4258 14912 4289
rect 14828 4252 14912 4258
rect 9984 3994 10432 4000
rect 17374 3873 17443 3874
rect 17502 3873 17569 3879
rect 17374 3867 17569 3873
rect 17374 3812 17508 3867
rect 17563 3812 17569 3867
rect 14877 3805 15139 3811
rect 14877 3746 15010 3805
rect 15069 3746 15139 3805
rect 14877 3740 15139 3746
rect 17374 3806 17569 3812
rect 10817 3455 10944 3461
rect 10944 3328 11647 3455
rect 10817 3322 10944 3328
rect 3732 3040 12000 3232
rect 14877 2950 14948 3740
rect 17374 2950 17443 3806
rect 17502 3800 17569 3806
rect 10817 2944 10944 2950
rect 14852 2830 18668 2950
rect 10817 2811 10944 2817
rect 992 -3736 1184 -2912
rect 800 -3928 1184 -3736
rect -8221 -6953 -7651 -6941
rect -8221 -7511 -8215 -6953
rect -7657 -7511 -7651 -6953
rect -8221 -7779 -7651 -7511
rect -8227 -8349 -8221 -7779
rect -7651 -8349 -7645 -7779
rect 18548 -8195 18668 2830
rect 18548 -8316 20035 -8195
rect 20156 -8316 20162 -8195
rect -15740 -10812 -13892 -10692
rect -14012 -12228 -13892 -10812
rect 18548 -12228 18668 -8316
rect -14012 -12348 18668 -12228
rect 18548 -12406 18668 -12348
<< via1 >>
rect -4956 11748 -4388 12316
rect 16292 11748 16860 12316
rect 9984 4000 10432 4448
rect 18076 4446 18148 4452
rect 18076 4392 18082 4446
rect 18082 4392 18142 4446
rect 18142 4392 18148 4446
rect 10817 3328 10944 3455
rect 10817 2817 10944 2944
rect -8221 -8349 -7651 -7779
rect 20035 -8316 20156 -8195
<< metal2 >>
rect -4956 13017 -4388 13022
rect -4960 12395 -4951 13017
rect -4393 12395 -4384 13017
rect 16292 13015 16860 13020
rect -4956 12316 -4388 12395
rect 16288 12393 16297 13015
rect 16855 12393 16864 13015
rect -4956 11742 -4388 11748
rect 16292 12316 16860 12393
rect 16292 11742 16860 11748
rect 13441 4865 20799 4992
rect 9978 4000 9984 4448
rect 10432 4000 10438 4448
rect 9984 3936 10432 4000
rect -15168 544 -3488 608
rect -15168 448 -15040 544
rect -3552 288 -3488 544
rect 2784 288 2848 3700
rect 9975 3488 9984 3936
rect 10432 3488 10441 3936
rect 10811 3328 10817 3455
rect 10944 3328 10950 3455
rect 10817 2944 10944 3328
rect 13441 2944 13568 4865
rect 18082 4452 18142 4865
rect 18070 4392 18076 4452
rect 18148 4392 18154 4452
rect 20672 3968 20799 4865
rect 20672 3832 20799 3841
rect 10811 2817 10817 2944
rect 10944 2817 13568 2944
rect -3552 224 2848 288
rect -8221 -7779 -7651 -7773
rect 20035 -8195 20156 -8189
rect 20156 -8316 20291 -8195
rect 20412 -8316 20421 -8195
rect 20035 -8322 20156 -8316
rect -8221 -8744 -7651 -8349
rect -8225 -9304 -8216 -8744
rect -7656 -9304 -7647 -8744
rect -8221 -9309 -7651 -9304
<< via2 >>
rect -4951 12395 -4393 13017
rect 16297 12393 16855 13015
rect 9984 3488 10432 3936
rect 20672 3841 20799 3968
rect 20291 -8316 20412 -8195
rect -8216 -9304 -7656 -8744
<< metal3 >>
rect -15808 13017 25984 13500
rect -15808 12395 -4951 13017
rect -4393 13015 25984 13017
rect -4393 12395 16297 13015
rect -15808 12393 16297 12395
rect 16855 12831 25984 13015
rect 16855 12513 24941 12831
rect 25259 12513 25984 12831
rect 16855 12393 25984 12513
rect -15808 12390 25984 12393
rect -4160 12388 25984 12390
rect 19496 4608 19672 12388
rect 15872 4480 19672 4608
rect 5539 3936 9821 3997
rect 15872 3968 16000 4480
rect 18344 4432 19672 4480
rect 9979 3936 10437 3941
rect 5539 3488 9984 3936
rect 10432 3488 10437 3936
rect 5539 3427 9821 3488
rect 9979 3483 10437 3488
rect -8221 -8744 -7651 -8739
rect -8221 -9304 -8216 -8744
rect -7656 -9304 -7651 -8744
rect -8221 -12771 -7651 -9304
rect 5539 -12771 6109 3427
rect 15360 3136 15488 3520
rect 17804 3184 17980 4024
rect 18344 3704 18520 4432
rect 20667 3968 20804 3973
rect 20667 3841 20672 3968
rect 20799 3841 20804 3968
rect 20667 3836 20804 3841
rect 17804 3136 19288 3184
rect 15360 3008 19288 3136
rect 19112 -12771 19288 3008
rect 20483 -8125 20796 -8004
rect 20286 -8194 20417 -8190
rect 20483 -8194 20604 -8125
rect 20286 -8195 20604 -8194
rect 20286 -8316 20291 -8195
rect 20412 -8315 20604 -8195
rect 20412 -8316 20417 -8315
rect 20286 -8321 20417 -8316
rect 25600 -12289 25920 -12288
rect 25595 -12607 25601 -12289
rect 25919 -12607 25925 -12289
rect 25600 -12771 25920 -12607
rect -15837 -14109 25949 -12771
<< via3 >>
rect 24941 12513 25259 12831
rect 25601 -12607 25919 -12289
<< metal4 >>
rect 24940 12831 25260 12832
rect 24940 12513 24941 12831
rect 25259 12513 25260 12831
rect 24940 7456 25260 12513
rect 25600 -12289 25920 -11232
rect 25600 -12607 25601 -12289
rect 25919 -12607 25920 -12289
rect 25600 -12608 25920 -12607
use JNW_VIS_ITIME  x1 ../JNW_GR02_SKY130A
timestamp 1744542523
transform 1 0 9649 0 1 12525
box -4353 -24590 9980 -1992
use JNW_VIS_TI  x2 ../JNW_GR02_SKY130A
timestamp 1744543763
transform 1 0 -5504 0 1 13448
box -9344 -19400 9900 -2398
use JNWTR_DFTSPCX1_CV  x3 ../JNW_TR_SKY130A
timestamp 1744542523
transform 1 0 14690 0 1 3314
box -150 -120 2130 1080
use JNWTR_DFTSPCX1_CV  x4
timestamp 1744542523
transform 1 0 17174 0 1 3320
box -150 -120 2130 1080
use dig  x5 ../JNW_GR02_SKY130A
timestamp 1744553953
transform 1 0 20732 0 1 -13844
box 0 1368 6600 22432
<< labels >>
flabel metal3 -15836 12390 -4951 12958 0 FreeSans 1600 0 0 0 VDD_1V8
port 0 nsew
flabel metal3 -15168 448 -15040 576 0 FreeSans 1600 0 0 0 PWR_UP_1V8
port 11 nsew
flabel space 27272 -12476 27332 -12356 0 FreeSans 1600 0 0 0 I_TEMP_OUT0
port 19 nsew
flabel space 27272 -9484 27332 -9364 0 FreeSans 1600 0 0 0 I_TEMP_OUT1
port 18 nsew
flabel space 27272 -6492 27332 -6372 0 FreeSans 1600 0 0 0 I_TEMP_OUT2
port 17 nsew
flabel space 27272 -3500 27332 -3380 0 FreeSans 1600 0 0 0 I_TEMP_OUT3
port 16 nsew
flabel space 27272 -508 27332 -388 0 FreeSans 1600 0 0 0 I_TEMP_OUT4
port 15 nsew
flabel space 27272 2484 27332 2604 0 FreeSans 1600 0 0 0 I_TEMP_OUT5
port 14 nsew
flabel space 27272 5476 27332 5596 0 FreeSans 1600 0 0 0 I_TEMP_OUT6
port 13 nsew
flabel space 27272 8468 27332 8588 0 FreeSans 1600 0 0 0 I_TEMP_OUT7
port 12 nsew
flabel metal3 -15808 -13312 -15104 -13120 0 FreeSans 1600 0 0 0 VSS
port 1 nsew
flabel metal3 -15740 -10812 -13892 -10692 0 FreeSans 1600 0 0 0 CLK
port 21 nsew
<< properties >>
string FIXED_BBOX 0 0 22267 11539
<< end >>
