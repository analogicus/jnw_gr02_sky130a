magic
tech sky130A
magscale 1 2
timestamp 1744379089
<< locali >>
rect 524 -2410 9684 -2404
rect 524 -2590 1678 -2410
rect 1858 -2590 3478 -2410
rect 3658 -2590 5278 -2410
rect 5458 -2590 7078 -2410
rect 7258 -2590 8858 -2410
rect 9038 -2590 9684 -2410
rect 524 -2596 9684 -2590
rect 524 -8044 716 -2596
rect 1288 -3824 1480 -2596
rect 2312 -3824 2504 -2596
rect 3088 -2824 3280 -2596
rect 4240 -2824 4432 -2596
rect 4888 -2836 5080 -2596
rect 6040 -2836 6232 -2596
rect 6688 -2836 6880 -2596
rect 7840 -2824 8032 -2596
rect 8468 -4424 8660 -2596
rect 9492 -4424 9684 -2596
rect 2000 -5280 2620 -5040
rect 3088 -5656 3464 -5464
rect 3644 -5656 4432 -5464
rect 3088 -5824 3280 -5656
rect 4240 -5824 4432 -5656
rect 4888 -5636 5284 -5444
rect 5476 -5636 6232 -5444
rect 4888 -5824 5080 -5636
rect 6040 -5836 6232 -5636
rect 6688 -5636 7064 -5444
rect 7256 -5636 8032 -5444
rect 6688 -5824 6880 -5636
rect 7840 -5824 8032 -5636
rect 8468 -5636 8844 -5444
rect 9036 -5636 9816 -5444
rect 8468 -5824 8660 -5636
rect 9624 -5816 9816 -5636
rect -9344 -8236 716 -8044
rect -9344 -13644 -9152 -8236
rect 1216 -8691 1328 -8072
rect 2084 -8184 2632 -8072
rect 931 -8915 5089 -8691
rect 931 -9787 1189 -8915
rect 2084 -9787 2581 -8915
rect 3504 -9787 4001 -9786
rect 4876 -9787 5089 -8915
rect 931 -10284 5089 -9787
rect 931 -11187 1189 -10284
rect 2084 -11139 2581 -10284
rect 3504 -11139 4001 -10284
rect 4876 -11139 5089 -10284
rect 6168 -10044 6360 -9820
rect 7832 -10044 8024 -9820
rect 6168 -10050 8024 -10044
rect 6168 -10230 6558 -10050
rect 6738 -10230 8024 -10050
rect 6168 -10236 8024 -10230
rect 6168 -11139 6360 -10236
rect 2036 -11187 6362 -11139
rect 931 -11684 6362 -11187
rect 931 -12472 1189 -11684
rect -7256 -12584 -1244 -12472
rect -80 -12584 1189 -12472
rect 931 -12586 1189 -12584
rect 2084 -12586 2581 -11684
rect 3504 -12586 4001 -11684
rect 4876 -12584 5089 -11684
rect 4784 -12586 7096 -12584
rect 931 -12776 7096 -12586
rect 931 -12779 5089 -12776
rect 931 -12786 1189 -12779
rect -9344 -13836 -7544 -13644
rect 6904 -18584 7096 -12776
rect 3984 -18636 7096 -18584
rect 3984 -18676 6156 -18636
rect 3984 -18764 5576 -18676
rect 5664 -18724 6156 -18676
rect 6244 -18724 7096 -18636
rect 5664 -18764 7096 -18724
rect 3984 -18776 7096 -18764
<< viali >>
rect 1678 -2590 1858 -2410
rect 3478 -2590 3658 -2410
rect 5278 -2590 5458 -2410
rect 7078 -2590 7258 -2410
rect 8858 -2590 9038 -2410
rect 1610 -5250 1790 -5070
rect 3464 -5656 3644 -5464
rect 5284 -5636 5476 -5444
rect 7064 -5636 7256 -5444
rect 8844 -5636 9036 -5444
rect -8590 -9630 -8410 -9450
rect -7740 -9680 -7500 -9440
rect -6434 -9674 -6206 -9446
rect -5956 -9668 -5716 -9440
rect -4636 -9680 -4396 -9452
rect -4156 -9668 -3916 -9440
rect -2836 -9680 -2596 -9452
rect -2356 -9668 -2116 -9440
rect -1036 -9680 -796 -9452
rect -597 -9697 -322 -9422
rect 6558 -10230 6738 -10050
rect 6156 -18724 6244 -18636
<< metal1 >>
rect 1672 -2410 1864 -2398
rect 1672 -2590 1678 -2410
rect 1858 -2590 1864 -2410
rect 1672 -4036 1864 -2590
rect 3472 -2410 3664 -2398
rect 3472 -2590 3478 -2410
rect 3658 -2590 3664 -2410
rect 3472 -3056 3664 -2590
rect 5272 -2410 5464 -2398
rect 5272 -2590 5278 -2410
rect 5458 -2590 5464 -2410
rect 5272 -3036 5464 -2590
rect 7072 -2410 7264 -2398
rect 7072 -2590 7078 -2410
rect 7258 -2590 7264 -2410
rect 7072 -2976 7264 -2590
rect 8852 -2410 9044 -2398
rect 8852 -2590 8858 -2410
rect 9038 -2590 9044 -2410
rect 1544 -4524 1608 -4348
rect 1928 -4524 2120 -4184
rect 3344 -4452 3408 -3288
rect 1544 -4668 2120 -4524
rect 3472 -4636 3664 -3144
rect 3856 -4616 4048 -3204
rect 5144 -4492 5208 -3288
rect 5272 -4636 5464 -3204
rect 5656 -4626 5848 -3204
rect 6944 -4452 7008 -3328
rect 7072 -4656 7264 -3204
rect 7456 -4616 7648 -3144
rect 8852 -4656 9044 -2590
rect 1544 -4724 2772 -4668
rect 1604 -4732 2772 -4724
rect 1604 -5070 1796 -4732
rect 1604 -5250 1610 -5070
rect 1790 -5250 1796 -5070
rect 1604 -5262 1796 -5250
rect 2708 -5388 2772 -4732
rect 3344 -5188 3408 -4968
rect 3856 -5144 4048 -4784
rect 3344 -5258 3408 -5252
rect 3464 -5336 4048 -5144
rect 5144 -5200 5208 -4968
rect 5656 -5200 5848 -4784
rect 5144 -5258 5208 -5252
rect 5284 -5336 5848 -5200
rect 6944 -5188 7008 -4968
rect 7456 -5124 7648 -4804
rect 6944 -5258 7008 -5252
rect 7064 -5316 7648 -5124
rect 8221 -5181 8300 -5175
rect 8724 -5188 8788 -4968
rect 9108 -5124 9300 -4784
rect 8724 -5258 8788 -5252
rect 3264 -5388 3424 -5376
rect 2708 -5452 3348 -5388
rect 3412 -5452 3424 -5388
rect 3464 -5452 3656 -5336
rect 3264 -5464 3424 -5452
rect 3458 -5464 3656 -5452
rect 3344 -5776 3408 -5464
rect 3458 -5656 3464 -5464
rect 3644 -5656 3656 -5464
rect 3458 -5668 3656 -5656
rect 3464 -6016 3656 -5668
rect 5144 -5388 5208 -5382
rect 5284 -5438 5476 -5336
rect 6944 -5388 7008 -5382
rect 5144 -5776 5208 -5452
rect 5278 -5444 5482 -5438
rect 5278 -5636 5284 -5444
rect 5476 -5636 5482 -5444
rect 5278 -5642 5482 -5636
rect 7064 -5438 7256 -5316
rect 5284 -5936 5476 -5642
rect 6944 -5776 7008 -5452
rect 7058 -5444 7262 -5438
rect 7058 -5636 7064 -5444
rect 7256 -5636 7262 -5444
rect 7058 -5642 7262 -5636
rect 7064 -5976 7256 -5642
rect 8221 -5712 8300 -5260
rect 8844 -5316 9300 -5124
rect 8724 -5388 8788 -5382
rect 8844 -5438 9036 -5316
rect 7456 -5904 8356 -5712
rect 8724 -5776 8788 -5452
rect 8838 -5444 9042 -5438
rect 8838 -5636 8844 -5444
rect 9036 -5636 9042 -5444
rect 8838 -5642 9042 -5636
rect 8844 -6036 9036 -5642
rect 3344 -7392 3408 -6288
rect 3472 -7636 3664 -6164
rect 3856 -7636 4048 -6144
rect 5144 -7412 5208 -6328
rect 5272 -7616 5464 -6164
rect 5656 -7616 5848 -6184
rect 6944 -7392 7008 -6348
rect 7072 -7656 7264 -6244
rect 7456 -7596 7648 -6204
rect 8724 -7412 8788 -6308
rect 8852 -7636 9044 -6184
rect 9236 -7556 9428 -6184
rect 3856 -8364 4048 -7784
rect -8596 -8556 4048 -8364
rect -8596 -9450 -8404 -8556
rect -5956 -9380 -320 -9140
rect -8596 -9630 -8590 -9450
rect -8410 -9630 -8404 -9450
rect -8596 -9642 -8404 -9630
rect -7791 -9440 -7249 -9429
rect -5956 -9434 -5716 -9380
rect -4156 -9434 -3916 -9380
rect -2356 -9434 -2116 -9380
rect -560 -9416 -320 -9380
rect 237 -9416 4623 -9196
rect -609 -9422 4623 -9416
rect -5968 -9440 -5704 -9434
rect -7791 -9680 -7740 -9440
rect -7500 -9446 -6194 -9440
rect -7500 -9674 -6434 -9446
rect -6206 -9674 -6194 -9446
rect -5968 -9668 -5956 -9440
rect -5716 -9668 -5704 -9440
rect -4168 -9440 -3904 -9434
rect -5968 -9674 -5704 -9668
rect -4648 -9452 -4384 -9446
rect -7500 -9680 -6194 -9674
rect -4648 -9680 -4636 -9452
rect -4396 -9680 -4384 -9452
rect -4168 -9668 -4156 -9440
rect -3916 -9668 -3904 -9440
rect -2368 -9440 -2104 -9434
rect -4168 -9674 -3904 -9668
rect -2848 -9452 -2584 -9446
rect -7791 -9691 -7249 -9680
rect -7022 -12988 -6958 -9680
rect -6680 -9760 -6440 -9680
rect -4648 -9686 -4384 -9680
rect -2848 -9680 -2836 -9452
rect -2596 -9680 -2584 -9452
rect -2368 -9668 -2356 -9440
rect -2116 -9668 -2104 -9440
rect -2368 -9674 -2104 -9668
rect -1048 -9452 -784 -9446
rect -2848 -9686 -2584 -9680
rect -1048 -9680 -1036 -9452
rect -796 -9680 -784 -9452
rect -1048 -9686 -784 -9680
rect -4636 -9760 -4396 -9686
rect -2836 -9760 -2596 -9686
rect -1036 -9760 -796 -9686
rect -609 -9697 -597 -9422
rect -322 -9483 4623 -9422
rect -322 -9697 524 -9483
rect -609 -9703 524 -9697
rect -6680 -10000 -760 -9760
rect 1467 -12016 1754 -9483
rect 2944 -10664 3136 -10658
rect 2944 -10862 3136 -10856
rect 4336 -12016 4623 -9483
rect 5656 -10664 5848 -7804
rect 7456 -8676 7648 -7744
rect 6028 -8962 6488 -8898
rect 6028 -10348 6092 -8962
rect 6552 -9536 6744 -8764
rect 9236 -9096 9428 -7804
rect 6428 -9748 6492 -9742
rect 6428 -9818 6492 -9812
rect 6552 -10050 6744 -9668
rect 6552 -10230 6558 -10050
rect 6738 -10230 6744 -10050
rect 6552 -10242 6744 -10230
rect 7448 -10348 7640 -9704
rect 8358 -9748 8422 -9742
rect 8422 -9812 8552 -9748
rect 8358 -9818 8422 -9812
rect 6028 -10412 7640 -10348
rect 7448 -10584 7640 -10412
rect 5228 -10856 5234 -10664
rect 5426 -10856 5848 -10664
rect 6464 -10776 7640 -10584
rect 1467 -12303 4623 -12016
rect -7022 -13052 -1322 -12988
rect -1258 -13052 -1252 -12988
rect 1088 -13008 1152 -13002
rect 1152 -13072 2988 -13008
rect 3052 -13072 3058 -13008
rect 1088 -13078 1152 -13072
rect -1322 -14028 -1258 -14022
rect -1322 -15512 -1258 -14092
rect 1088 -14068 1152 -14062
rect 1088 -15512 1152 -14132
rect 6504 -16390 6696 -10776
rect 6504 -16490 6530 -16390
rect 6630 -16490 6696 -16390
rect 6504 -16556 6696 -16490
rect 5704 -17376 6504 -17184
rect 6144 -18470 6150 -18370
rect 6250 -18470 6256 -18370
rect 6150 -18636 6250 -18470
rect 6150 -18724 6156 -18636
rect 6244 -18724 6250 -18636
rect 6150 -18736 6250 -18724
<< via1 >>
rect 3344 -5252 3408 -5188
rect 5144 -5252 5208 -5200
rect 6944 -5252 7008 -5188
rect 8221 -5260 8300 -5181
rect 8724 -5252 8788 -5188
rect 3348 -5452 3412 -5388
rect 5144 -5452 5208 -5388
rect 6944 -5452 7008 -5388
rect 8724 -5452 8788 -5388
rect 2944 -10856 3136 -10664
rect 6428 -9812 6492 -9748
rect 8358 -9812 8422 -9748
rect 5234 -10856 5426 -10664
rect -1322 -13052 -1258 -12988
rect 1088 -13072 1152 -13008
rect 2988 -13072 3052 -13008
rect -1322 -14092 -1258 -14028
rect 1088 -14132 1152 -14068
rect 6530 -16490 6630 -16390
rect 6150 -18470 6250 -18370
<< metal2 >>
rect 8215 -5188 8221 -5181
rect 3338 -5252 3344 -5188
rect 3408 -5200 6944 -5188
rect 3408 -5252 5144 -5200
rect 5208 -5252 6944 -5200
rect 7008 -5252 8221 -5188
rect 8215 -5260 8221 -5252
rect 8300 -5188 8306 -5181
rect 8300 -5252 8724 -5188
rect 8788 -5252 8794 -5188
rect 8300 -5260 8306 -5252
rect 3342 -5452 3348 -5388
rect 3412 -5452 5144 -5388
rect 5208 -5452 6944 -5388
rect 7008 -5452 8724 -5388
rect 8788 -5452 8794 -5388
rect 6422 -9812 6428 -9748
rect 6492 -9812 8358 -9748
rect 8422 -9812 8428 -9748
rect 5234 -10664 5426 -10658
rect 2938 -10856 2944 -10664
rect 3136 -10856 5234 -10664
rect -1322 -12988 -1258 -12982
rect 2988 -13008 3052 -10856
rect 5234 -10862 5426 -10856
rect -1322 -14028 -1258 -13052
rect 1082 -13072 1088 -13008
rect 1152 -13072 1158 -13008
rect -1328 -14092 -1322 -14028
rect -1258 -14092 -1252 -14028
rect 1088 -14068 1152 -13072
rect 2988 -13078 3052 -13072
rect 1082 -14132 1088 -14068
rect 1152 -14132 1158 -14068
rect 6315 -16390 6405 -16386
rect 6310 -16395 6530 -16390
rect 6310 -16485 6315 -16395
rect 6405 -16485 6530 -16395
rect 6310 -16490 6530 -16485
rect 6630 -16490 6636 -16390
rect 6315 -16494 6405 -16490
rect 6150 -18215 6250 -18210
rect 6146 -18305 6155 -18215
rect 6245 -18305 6254 -18215
rect 6150 -18370 6250 -18305
rect 6150 -18476 6250 -18470
<< via2 >>
rect 6315 -16485 6405 -16395
rect 6155 -18305 6245 -18215
<< metal3 >>
rect 1270 -16390 1370 -16070
rect 4070 -16390 4170 -16070
rect 1250 -16490 3510 -16390
rect 3990 -16490 4170 -16390
rect 4370 -16395 6410 -16390
rect 4370 -16485 6315 -16395
rect 6405 -16485 6410 -16395
rect 4370 -16490 6410 -16485
rect 6150 -18071 6250 -18070
rect 6145 -18169 6151 -18071
rect 6249 -18169 6255 -18071
rect 6150 -18215 6250 -18169
rect 6150 -18305 6155 -18215
rect 6245 -18305 6250 -18215
rect 6150 -18310 6250 -18305
<< via3 >>
rect 6151 -18169 6249 -18071
<< metal4 >>
rect 1280 -16390 1380 -16080
rect 4180 -16390 4280 -16050
rect 5460 -16160 6250 -16060
rect 1130 -16490 4670 -16390
rect 6150 -18071 6250 -16160
rect 6150 -18169 6151 -18071
rect 6249 -18169 6250 -18071
rect 6150 -18170 6250 -18169
use JNWATR_NCH_12C5F0  JNWATR_NCH_12C5F0_0 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 6264 0 1 -9172
box -184 -128 1848 928
use JNWATR_NCH_12C5F0  JNWATR_NCH_12C5F0_1
timestamp 1734044400
transform 1 0 6264 0 1 -9972
box -184 -128 1848 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_0 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 6784 0 1 -3472
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_1
timestamp 1734044400
transform 1 0 6784 0 1 -4272
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_2
timestamp 1734044400
transform 1 0 6784 0 1 -5072
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_6
timestamp 1734044400
transform 1 0 3184 0 1 -3472
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_7
timestamp 1734044400
transform 1 0 3184 0 1 -4272
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_8
timestamp 1734044400
transform 1 0 3184 0 1 -5072
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_9
timestamp 1734044400
transform 1 0 4984 0 1 -5072
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_10
timestamp 1734044400
transform 1 0 4984 0 1 -4272
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_11
timestamp 1734044400
transform 1 0 4984 0 1 -3472
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_16
timestamp 1734044400
transform 1 0 8564 0 1 -8072
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_17
timestamp 1734044400
transform 1 0 8564 0 1 -7272
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_18
timestamp 1734044400
transform 1 0 3184 0 1 -6472
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_21
timestamp 1734044400
transform 1 0 6784 0 1 -6472
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_22
timestamp 1734044400
transform 1 0 6784 0 1 -8072
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_23
timestamp 1734044400
transform 1 0 6784 0 1 -7272
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_24
timestamp 1734044400
transform 1 0 4984 0 1 -6472
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_25
timestamp 1734044400
transform 1 0 3184 0 1 -8072
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_26
timestamp 1734044400
transform 1 0 3184 0 1 -7272
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_27
timestamp 1734044400
transform 1 0 8564 0 1 -6472
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_28
timestamp 1734044400
transform 1 0 4984 0 1 -8072
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_29
timestamp 1734044400
transform 1 0 4984 0 1 -7272
box -184 -128 1336 928
use JNWTR_CAPX4  JNWTR_CAPX4_0 ../JNW_TR_SKY130A
timestamp 1744372914
transform -1 0 6030 0 -1 -16390
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_1
timestamp 1744372914
transform 1 0 -430 0 1 -16160
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_2
timestamp 1744372914
transform -1 0 3160 0 -1 -16390
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_3
timestamp 1744372914
transform 1 0 2440 0 1 -16160
box 480 0 3120 2640
use JNWTR_RPPO2  JNWTR_RPPO2_0 ../JNW_TR_SKY130A
timestamp 1744291457
transform -1 0 48 0 1 -12600
box 0 0 1448 3440
use JNWTR_RPPO2  JNWTR_RPPO2_1
timestamp 1744291457
transform -1 0 -5352 0 1 -12600
box 0 0 1448 3440
use JNWTR_RPPO2  JNWTR_RPPO2_2
timestamp 1744291457
transform -1 0 -3552 0 1 -12600
box 0 0 1448 3440
use JNWTR_RPPO2  JNWTR_RPPO2_3
timestamp 1744291457
transform -1 0 -1752 0 1 -12600
box 0 0 1448 3440
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1734020192
transform 1 0 980 0 1 -11400
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1734020192
transform 1 0 2380 0 1 -11400
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1734020192
transform 1 0 3780 0 1 -11400
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1734020192
transform 1 0 3780 0 1 -10000
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1734020192
transform 1 0 980 0 1 -10000
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1734020192
transform 1 0 3780 0 1 -12800
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1734020192
transform 1 0 980 0 1 -12800
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8
timestamp 1734020192
transform 1 0 2380 0 1 -12800
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_9
timestamp 1734020192
transform 1 0 2380 0 1 -10000
box 0 0 1340 1340
use JNWATR_PCH_2C5F0  x2 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 8564 0 1 -5072
box -184 -128 1208 928
use JNWTR_RPPO2  x3
timestamp 1744291457
transform -1 0 2648 0 1 -8200
box 0 0 1448 3440
use JNW_VIS_OTA  x7 ../JNW_GR02_SKY130A
timestamp 1744372914
transform 1 0 1120 0 1 -16000
box -9120 -3400 4936 2656
use JNWTR_RPPO4  x14 ../JNW_TR_SKY130A
timestamp 1744372914
transform -1 0 -7120 0 1 -12600
box 0 0 1880 3440
use JNWATR_PCH_2C5F0  x15
timestamp 1734044400
transform 1 0 1384 0 1 -4472
box -184 -128 1208 928
<< labels >>
flabel metal1 -8596 -8556 -8404 -8364 0 FreeSans 1600 0 0 0 VREF
port 3 nsew
flabel metal1 9236 -9096 9428 -8904 0 FreeSans 1600 0 0 0 I_TEMP
port 4 nsew
flabel locali -9344 -8236 -9152 -8044 0 FreeSans 1600 0 0 0 VDD
port 5 nsew
flabel locali 6904 -18776 7096 -18584 0 FreeSans 1600 0 0 0 VSS
port 6 nsew
flabel metal1 6304 -17376 6496 -17184 0 FreeSans 1600 0 0 0 LPO
port 7 nsew
flabel metal1 6504 -15896 6696 -15704 0 FreeSans 1600 0 0 0 LPI
port 8 nsew
flabel metal1 8488 -9812 8552 -9748 0 FreeSans 1600 0 0 0 PWR_UP
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 2904 10680
<< end >>
