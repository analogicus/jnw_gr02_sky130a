** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_GR02_SKY130A/TB_JNW_VIS_TI.sch
**.subckt TB_JNW_VIS_TI VDD VSS VREF I_TEMP PWR_UP LPI LPO
*.ipin VDD
*.ipin VSS
*.opin VREF
*.opin I_TEMP
*.ipin PWR_UP
*.opin LPI
*.opin LPO
x1 VDD VREF LPI LPO I_TEMP PWR_UP VSS JNW_VIS_TI
**** begin user architecture code



.param mc_mm_switch=0
.param mc_pr_switch=0
.include tt.spi
*.include ss.spi
.option gmin=1e-15
.lib ../../../tech/ngspice/temperature.spi Tl
.lib ../../../tech/ngspice/supply.spi Vl
.include ../../../../cpdk/ngspice/ideal_circuits.spi
.include /home/domen/pro/aicex/ip/cpdk/ngspice/tian_subckt.lib

X999 LPI LPO loopgainprobe

VSS  VSS  0     dc 0
VDD  VDD VSS dc 1.8
VPUP PWR_UP VSS PULSE ( 0 1.8 1NS 1PS 1PS 1NS 1S 1)
VSENS I_TEMP 0 dc 0.5


.option temp = 25
.option savecurrents
.save all
.control

.IC V(LPO)=0.5
optran 0 0 0 10n 10u 0
op
write TB_JNW_VIS_TI.raw
exit
.endc
.end



**** end user architecture code
**.ends

* expanding   symbol:  JNW_GR02_SKY130A/JNW_VIS_TI.sym # of pins=7
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_GR02_SKY130A/JNW_VIS_TI.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_GR02_SKY130A/JNW_VIS_TI.sch
.subckt JNW_VIS_TI VDD VREF LPI LPO I_TEMP PWR_UP VSS
*.ipin VDD
*.ipin VSS
*.opin VREF
*.opin I_TEMP
*.ipin PWR_UP
*.opin LPI
*.opin LPO
XQ1 VSS VSS VIN sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1 mult=1
XQ2 VSS VSS VD2 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=8 mult=8
x7 VDD VIN VIP VSS LPO JNW_VIS_OTA
x11 VDD PWR_UP LPI VSS JNWATR_NCH_12C1F2
x1<0> LPI VSS JNWTR_CAPX1
x1<1> LPI VSS JNWTR_CAPX1
x1<2> LPI VSS JNWTR_CAPX1
x5<0> VIP VREF VSS JNWTR_RPPO8
x5<1> VIP VREF VSS JNWTR_RPPO8
x8<0> VD2 VIP VSS JNWTR_RPPO4
x8<1> VD2 VIP VSS JNWTR_RPPO4
x8<2> VD2 VIP VSS JNWTR_RPPO4
x8<3> VD2 VIP VSS JNWTR_RPPO4
x8<4> VD2 VIP VSS JNWTR_RPPO4
x8<5> VD2 VIP VSS JNWTR_RPPO4
x8<6> VD2 VIP VSS JNWTR_RPPO4
x1 net1 net1 VDD VDD JNWATR_PCH_8C1F2
x2 VIN net1 VDD VDD JNWATR_PCH_8C1F2
x3 VREF net1 VDD VDD JNWATR_PCH_8C1F2
x4 I_TEMP net1 VDD VDD JNWATR_PCH_8C1F2
x6 net1 LPI VSS VSS JNWATR_NCH_8C5F0
x2<0> VCAP VSS JNWTR_CAPX1
x2<1> VCAP VSS JNWTR_CAPX1
x2<2> VCAP VSS JNWTR_CAPX1
x2<3> VCAP VSS JNWTR_CAPX1
x2<4> VCAP VSS JNWTR_CAPX1
x2<5> VCAP VSS JNWTR_CAPX1
x2<6> VCAP VSS JNWTR_CAPX1
x2<7> VCAP VSS JNWTR_CAPX1
x2<8> VCAP VSS JNWTR_CAPX1
x2<9> VCAP VSS JNWTR_CAPX1
x2<10> VCAP VSS JNWTR_CAPX1
x2<11> VCAP VSS JNWTR_CAPX1
x2<12> VCAP VSS JNWTR_CAPX1
x2<13> VCAP VSS JNWTR_CAPX1
x2<14> VCAP VSS JNWTR_CAPX1
x2<15> VCAP VSS JNWTR_CAPX1
x2<16> VCAP VSS JNWTR_CAPX1
x2<17> VCAP VSS JNWTR_CAPX1
x2<18> VCAP VSS JNWTR_CAPX1
x2<19> VCAP VSS JNWTR_CAPX1
x2<20> VCAP VSS JNWTR_CAPX1
x2<21> VCAP VSS JNWTR_CAPX1
x2<22> VCAP VSS JNWTR_CAPX1
x2<23> VCAP VSS JNWTR_CAPX1
x2<24> VCAP VSS JNWTR_CAPX1
x2<25> VCAP VSS JNWTR_CAPX1
x2<26> VCAP VSS JNWTR_CAPX1
x2<27> VCAP VSS JNWTR_CAPX1
x2<28> VCAP VSS JNWTR_CAPX1
x2<29> VCAP VSS JNWTR_CAPX1
x2<30> VCAP VSS JNWTR_CAPX1
x2<31> VCAP VSS JNWTR_CAPX1
x2<32> VCAP VSS JNWTR_CAPX1
x2<33> VCAP VSS JNWTR_CAPX1
x2<34> VCAP VSS JNWTR_CAPX1
x2<35> VCAP VSS JNWTR_CAPX1
x2<36> VCAP VSS JNWTR_CAPX1
x2<37> VCAP VSS JNWTR_CAPX1
x2<38> VCAP VSS JNWTR_CAPX1
x2<39> VCAP VSS JNWTR_CAPX1
x2<40> VCAP VSS JNWTR_CAPX1
x2<41> VCAP VSS JNWTR_CAPX1
x2<42> VCAP VSS JNWTR_CAPX1
x2<43> VCAP VSS JNWTR_CAPX1
x2<44> VCAP VSS JNWTR_CAPX1
x2<45> VCAP VSS JNWTR_CAPX1
x2<46> VCAP VSS JNWTR_CAPX1
x2<47> VCAP VSS JNWTR_CAPX1
x2<48> VCAP VSS JNWTR_CAPX1
x2<49> VCAP VSS JNWTR_CAPX1
x2<50> VCAP VSS JNWTR_CAPX1
x2<51> VCAP VSS JNWTR_CAPX1
x2<52> VCAP VSS JNWTR_CAPX1
x2<53> VCAP VSS JNWTR_CAPX1
x2<54> VCAP VSS JNWTR_CAPX1
x2<55> VCAP VSS JNWTR_CAPX1
x2<56> VCAP VSS JNWTR_CAPX1
x2<57> VCAP VSS JNWTR_CAPX1
x2<58> VCAP VSS JNWTR_CAPX1
x2<59> VCAP VSS JNWTR_CAPX1
x2<60> VCAP VSS JNWTR_CAPX1
x2<61> VCAP VSS JNWTR_CAPX1
x2<62> VCAP VSS JNWTR_CAPX1
x2<63> VCAP VSS JNWTR_CAPX1
x2<64> VCAP VSS JNWTR_CAPX1
x2<65> VCAP VSS JNWTR_CAPX1
x2<66> VCAP VSS JNWTR_CAPX1
x2<67> VCAP VSS JNWTR_CAPX1
x2<68> VCAP VSS JNWTR_CAPX1
x2<69> VCAP VSS JNWTR_CAPX1
x2<70> VCAP VSS JNWTR_CAPX1
x2<71> VCAP VSS JNWTR_CAPX1
x2<72> VCAP VSS JNWTR_CAPX1
x2<73> VCAP VSS JNWTR_CAPX1
x2<74> VCAP VSS JNWTR_CAPX1
x2<75> VCAP VSS JNWTR_CAPX1
x2<76> VCAP VSS JNWTR_CAPX1
x2<77> VCAP VSS JNWTR_CAPX1
x2<78> VCAP VSS JNWTR_CAPX1
x2<79> VCAP VSS JNWTR_CAPX1
x2<80> VCAP VSS JNWTR_CAPX1
x2<81> VCAP VSS JNWTR_CAPX1
x2<82> VCAP VSS JNWTR_CAPX1
x2<83> VCAP VSS JNWTR_CAPX1
x2<84> VCAP VSS JNWTR_CAPX1
x2<85> VCAP VSS JNWTR_CAPX1
x2<86> VCAP VSS JNWTR_CAPX1
x2<87> VCAP VSS JNWTR_CAPX1
x2<88> VCAP VSS JNWTR_CAPX1
x2<89> VCAP VSS JNWTR_CAPX1
x2<90> VCAP VSS JNWTR_CAPX1
x2<91> VCAP VSS JNWTR_CAPX1
x2<92> VCAP VSS JNWTR_CAPX1
x2<93> VCAP VSS JNWTR_CAPX1
x2<94> VCAP VSS JNWTR_CAPX1
x2<95> VCAP VSS JNWTR_CAPX1
x2<96> VCAP VSS JNWTR_CAPX1
x2<97> VCAP VSS JNWTR_CAPX1
x2<98> VCAP VSS JNWTR_CAPX1
x2<99> VCAP VSS JNWTR_CAPX1
x2<100> VCAP VSS JNWTR_CAPX1
x5 VCAP net1 VDD VDD JNWATR_PCH_8C1F2
.ends


* expanding   symbol:  JNW_GR02_SKY130A/JNW_VIS_OTA.sym # of pins=5
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_GR02_SKY130A/JNW_VIS_OTA.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_GR02_SKY130A/JNW_VIS_OTA.sch
.subckt JNW_VIS_OTA VDD VIN VIP VSS VOUT
*.ipin VDD
*.ipin VIP
*.ipin VIN
*.ipin VSS
*.opin VOUT
x1 V2 VIP VOP VOP JNWATR_PCH_4C1F2
x10 V1 VIN VOP VOP JNWATR_PCH_4C1F2
x3 VOUT V1 VSS VSS JNWATR_NCH_4C5F0
x4 V2 V2 VSS VSS JNWATR_NCH_4C5F0
x5 net1 V2 VSS VSS JNWATR_NCH_4C5F0
x6 V1 V1 VSS VSS JNWATR_NCH_4C5F0
x7 VOUT net1 VDD VDD JNWATR_PCH_12C5F0
x8<0> VOP VGS_M VDD VDD JNWATR_PCH_8C1F2
x8<1> VOP VGS_M VDD VDD JNWATR_PCH_8C1F2
x9 VGS_M VGS_M VDD VDD JNWATR_PCH_8C1F2
x11 net1 net1 VDD VDD JNWATR_PCH_12C5F0
x2<0> VSS net2 VSS JNWTR_RPPO4
x1<0> net2 VGS_M VSS JNWTR_RPPO4
x1<1> net2 VGS_M VSS JNWTR_RPPO4
x1<2> net2 VGS_M VSS JNWTR_RPPO4
x1<3> net2 VGS_M VSS JNWTR_RPPO4
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_12C1F2.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_12C1F2.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_12C1F2.sch
.subckt JNWATR_NCH_12C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.22 W=8.32 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_CAPX1.sym # of pins=2
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sch
.subckt JNWTR_CAPX1 A B
*.iopin A
*.iopin B
XC1 B A sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RPPO8.sym # of pins=3
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO8.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO8.sch
.subckt JNWTR_RPPO8 N P B
*.iopin P
*.iopin N
*.iopin B
XXA1 N P B JNWTR_RES8
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RPPO4.sym # of pins=3
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO4.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO4.sch
.subckt JNWTR_RPPO4 N P B
*.iopin P
*.iopin N
*.iopin B
XXA1 N P B JNWTR_RES4
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_8C1F2.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_8C1F2.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_8C1F2.sch
.subckt JNWATR_PCH_8C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.22 W=5.76 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_8C5F0.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_8C5F0.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_8C5F0.sch
.subckt JNWATR_NCH_8C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.94 W=5.76 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_4C1F2.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C1F2.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C1F2.sch
.subckt JNWATR_PCH_4C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.22 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sch
.subckt JNWATR_NCH_4C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.94 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_12C5F0.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_12C5F0.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_12C5F0.sch
.subckt JNWATR_PCH_12C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.94 W=8.32 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RES8.sym # of pins=3
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RES8.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RES8.sch
.subckt JNWTR_RES8 N P B
*.iopin N
*.iopin P
*.iopin B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_1 INT_1 INT_0 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_2 INT_2 INT_1 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_3 INT_3 INT_2 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_4 INT_4 INT_3 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_5 INT_5 INT_4 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_6 INT_6 INT_5 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_7 P INT_6 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RES4.sym # of pins=3
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RES4.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RES4.sch
.subckt JNWTR_RES4 N P B
*.iopin N
*.iopin P
*.iopin B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_1 INT_1 INT_0 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_2 INT_2 INT_1 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_3 P INT_2 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
.ends

.end
