magic
tech sky130A
timestamp 1744131902
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_0 ~/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 -2408 0 1 2064
box -92 -64 924 464
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_1
timestamp 1734044400
transform 1 0 -3908 0 1 3364
box -92 -64 924 464
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_2
timestamp 1734044400
transform 1 0 -2408 0 1 2464
box -92 -64 924 464
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_3
timestamp 1734044400
transform 1 0 -2408 0 1 3264
box -92 -64 924 464
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_4
timestamp 1734044400
transform 1 0 -2408 0 1 2864
box -92 -64 924 464
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_5
timestamp 1734044400
transform 1 0 -3908 0 1 2164
box -92 -64 924 464
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_6
timestamp 1734044400
transform 1 0 -3908 0 1 2564
box -92 -64 924 464
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_7
timestamp 1734044400
transform 1 0 -3908 0 1 2964
box -92 -64 924 464
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_0 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 -3908 0 1 4764
box -92 -64 924 464
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_1
timestamp 1734044400
transform 1 0 -2408 0 -1 5164
box -92 -64 924 464
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_2
timestamp 1734044400
transform 1 0 -2408 0 1 5164
box -92 -64 924 464
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_3
timestamp 1734044400
transform 1 0 -2408 0 1 5564
box -92 -64 924 464
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_4
timestamp 1734044400
transform 1 0 -2408 0 1 5964
box -92 -64 924 464
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_5
timestamp 1734044400
transform 1 0 -3908 0 1 5964
box -92 -64 924 464
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_6
timestamp 1734044400
transform 1 0 -3908 0 1 5164
box -92 -64 924 464
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_7
timestamp 1734044400
transform 1 0 -3908 0 1 5564
box -92 -64 924 464
use JNWTR_RPPO2  JNWTR_RPPO2_0 ../JNW_TR_SKY130A
timestamp 1744131902
transform 1 0 2986 0 1 2001
box 0 0 724 1720
use JNWTR_RPPO2  JNWTR_RPPO2_1
timestamp 1744131902
transform 1 0 2000 0 1 4000
box 0 0 724 1720
use JNWTR_RPPO2  x6
timestamp 1744131902
transform 1 0 2000 0 1 2000
box 0 0 724 1720
use JNWATR_PCH_12C5F0  xa01
timestamp 1734044400
transform 1 0 -908 0 1 2064
box -92 -64 924 464
use JNWATR_PCH_12C5F0  xa02
timestamp 1734044400
transform 1 0 -908 0 1 2464
box -92 -64 924 464
use JNWATR_NCH_12C5F0  xc01 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 340 0 1 2020
box -92 -64 924 464
use JNWATR_NCH_12C5F0  xc02
timestamp 1734044400
transform 1 0 340 0 1 2420
box -92 -64 924 464
use JNWATR_NCH_12C5F0  xc03
timestamp 1734044400
transform 1 0 340 0 1 2820
box -92 -64 924 464
use JNWATR_NCH_12C5F0  xc04
timestamp 1734044400
transform 1 0 340 0 1 3220
box -92 -64 924 464
<< properties >>
string FIXED_BBOX 0 0 1172 3620
<< end >>
