magic
tech sky130A
magscale 1 2
timestamp 1744236000
<< checkpaint >>
rect 0 0 16424 3440
use JNWATR_NCH_12C5F0 x10 ../JNW_ATR_SKY130A
transform 1 0 0 0 1 0
box 0 0 1664 800
use JNWATR_PCH_12C5F0 x13 ../JNW_ATR_SKY130A
transform 1 0 1664 0 1 0
box 1664 0 3328 800
use JNWATR_PCH_12C5F0 x14 ../JNW_ATR_SKY130A
transform 1 0 3328 0 1 0
box 3328 0 4992 800
use JNWATR_PCH_12C1F2 x1_0 ../JNW_ATR_SKY130A
transform 1 0 4992 0 1 0
box 4992 0 6656 800
use JNWATR_PCH_12C1F2 x1_1 ../JNW_ATR_SKY130A
transform 1 0 4992 0 1 800
box 4992 800 6656 1600
use JNWATR_PCH_12C1F2 x1_2 ../JNW_ATR_SKY130A
transform 1 0 4992 0 1 1600
box 4992 1600 6656 2400
use JNWATR_PCH_12C1F2 x1_3 ../JNW_ATR_SKY130A
transform 1 0 4992 0 1 2400
box 4992 2400 6656 3200
use JNWATR_NCH_12C5F0 x2 ../JNW_ATR_SKY130A
transform 1 0 6656 0 1 0
box 6656 0 8320 800
use JNWATR_PCH_12C5F0 x2_0 ../JNW_ATR_SKY130A
transform 1 0 8320 0 1 0
box 8320 0 9984 800
use JNWATR_PCH_12C5F0 x2_1 ../JNW_ATR_SKY130A
transform 1 0 8320 0 1 800
box 8320 800 9984 1600
use JNWATR_PCH_12C5F0 x2_2 ../JNW_ATR_SKY130A
transform 1 0 8320 0 1 1600
box 8320 1600 9984 2400
use JNWATR_PCH_12C5F0 x2_3 ../JNW_ATR_SKY130A
transform 1 0 8320 0 1 2400
box 8320 2400 9984 3200
use JNWATR_NCH_12C5F0 x3 ../JNW_ATR_SKY130A
transform 1 0 9984 0 1 0
box 9984 0 11648 800
use JNWATR_PCH_12C5F0 x3_0 ../JNW_ATR_SKY130A
transform 1 0 11648 0 1 0
box 11648 0 13312 800
use JNWATR_PCH_12C5F0 x3_1 ../JNW_ATR_SKY130A
transform 1 0 11648 0 1 800
box 11648 800 13312 1600
use JNWATR_PCH_12C5F0 x3_2 ../JNW_ATR_SKY130A
transform 1 0 11648 0 1 1600
box 11648 1600 13312 2400
use JNWATR_PCH_12C5F0 x3_3 ../JNW_ATR_SKY130A
transform 1 0 11648 0 1 2400
box 11648 2400 13312 3200
use JNWATR_NCH_12C5F0 x5 ../JNW_ATR_SKY130A
transform 1 0 13312 0 1 0
box 13312 0 14976 800
use JNWTR_RPPO2 x6 ../JNW_TR_SKY130A
transform 1 0 14976 0 1 0
box 14976 0 16424 3440
use JNWATR_PCH_12C1F2 x7_0 ../JNW_ATR_SKY130A
transform 1 0 0 0 1 3440
box 0 3440 1664 4240
use JNWATR_PCH_12C1F2 x7_1 ../JNW_ATR_SKY130A
transform 1 0 0 0 1 4240
box 0 4240 1664 5040
use JNWATR_PCH_12C1F2 x7_2 ../JNW_ATR_SKY130A
transform 1 0 0 0 1 5040
box 0 5040 1664 5840
use JNWATR_PCH_12C1F2 x7_3 ../JNW_ATR_SKY130A
transform 1 0 0 0 1 5840
box 0 5840 1664 6640
use JNWTR_RPPO2 x8_0 ../JNW_TR_SKY130A
transform 1 0 1664 0 1 3440
box 1664 3440 3112 6880
use JNWTR_RPPO2 x8_1 ../JNW_TR_SKY130A
transform 1 0 1664 0 1 6880
box 1664 6880 3112 10320
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 16424 3440
<< end >>
