magic
tech sky130A
magscale 1 2
timestamp 1745488630
<< dnwell >>
rect 27800 -11000 33000 -200
<< nwell >>
rect 27400 -200 33400 200
rect 27400 -11000 27800 -200
rect 33000 -11000 33400 -200
rect 27400 -11400 33400 -11000
<< locali >>
rect 23804 -1010 37352 -1004
rect 23804 -1190 25078 -1010
rect 25258 -1190 37352 -1010
rect 23804 -1196 37352 -1190
rect 24688 -2224 24880 -1196
rect 26352 -2224 26544 -1196
rect 36456 -1458 36632 -1196
rect 29556 -1550 30906 -1490
rect 24688 -7250 24880 -4920
rect 26352 -5304 26544 -4872
rect 26096 -5496 26556 -5304
rect 26096 -5672 26288 -5496
rect 24688 -7430 24690 -7250
rect 24870 -7430 24880 -7250
rect 24688 -8644 24880 -7430
rect 26096 -8644 26288 -6884
rect 22220 -8836 26288 -8644
rect 24688 -10024 24880 -8836
rect 28576 -9260 28796 -1970
rect 29556 -2610 29616 -1550
rect 29016 -3130 29076 -2790
rect 30276 -3130 30336 -2810
rect 29016 -3142 30336 -3130
rect 29016 -3190 30276 -3142
rect 29556 -3970 29616 -3190
rect 29016 -4530 29076 -4230
rect 30276 -4530 30336 -4230
rect 29016 -4542 30336 -4530
rect 29016 -4590 30276 -4542
rect 29556 -5450 29616 -4590
rect 29016 -5970 29076 -5610
rect 30276 -5970 30336 -5630
rect 29016 -5982 30336 -5970
rect 29016 -6030 30276 -5982
rect 29556 -6870 29616 -6030
rect 29016 -7370 29076 -7030
rect 30276 -7370 30336 -7030
rect 29016 -7382 30336 -7370
rect 29016 -7430 30276 -7382
rect 29556 -8270 29616 -7430
rect 29016 -8770 29076 -8410
rect 30276 -8770 30336 -8410
rect 30576 -8720 30756 -1838
rect 30846 -5430 30906 -1550
rect 36456 -1622 36462 -1458
rect 36626 -1622 36632 -1458
rect 36456 -1628 36632 -1622
rect 36006 -2010 36216 -1950
rect 35180 -4898 35372 -2164
rect 36156 -2630 36216 -2010
rect 35616 -3250 35676 -2830
rect 36876 -3250 36936 -2810
rect 35616 -3310 36936 -3250
rect 36156 -3970 36216 -3310
rect 35616 -4490 35676 -4150
rect 36876 -4490 36936 -4170
rect 37160 -4436 37352 -1196
rect 35616 -4496 36936 -4490
rect 35616 -4544 36292 -4496
rect 36340 -4544 36936 -4496
rect 35616 -4550 36936 -4544
rect 35180 -5062 35194 -4898
rect 35358 -5062 35372 -4898
rect 30846 -5490 31598 -5430
rect 30846 -8770 30906 -5490
rect 29016 -8782 30906 -8770
rect 29016 -8830 30276 -8782
rect 30336 -8830 30906 -8782
rect 28576 -9390 28796 -9380
rect 35180 -10024 35372 -5062
rect 24688 -10216 35372 -10024
<< viali >>
rect 25078 -1190 25258 -1010
rect 24690 -7430 24870 -7250
rect 30576 -1838 30756 -1670
rect 30276 -3190 30336 -3142
rect 30276 -4590 30336 -4542
rect 30276 -6030 30336 -5982
rect 30276 -7430 30336 -7382
rect 36462 -1622 36626 -1458
rect 36292 -4544 36340 -4496
rect 35194 -5062 35358 -4898
rect 31598 -5490 31646 -5430
rect 30276 -8830 30336 -8782
rect 28576 -9380 28796 -9260
<< metal1 >>
rect 25072 -1010 25264 -998
rect 25072 -1190 25078 -1010
rect 25258 -1190 25264 -1010
rect 25072 -2356 25264 -1190
rect 36456 -1458 36632 -1446
rect 36456 -1622 36462 -1458
rect 36626 -1622 36632 -1458
rect 25968 -1670 30772 -1664
rect 25968 -1672 30576 -1670
rect 25968 -1848 29856 -1672
rect 30032 -1838 30576 -1672
rect 30756 -1838 30772 -1670
rect 36456 -1692 36632 -1622
rect 30032 -1848 30772 -1838
rect 25968 -1856 30772 -1848
rect 25968 -2316 26160 -1856
rect 36450 -1868 36456 -1692
rect 36632 -1868 36638 -1692
rect 24944 -3092 25008 -2708
rect 25072 -3176 25264 -2408
rect 30264 -3142 30348 -3136
rect 30264 -3190 30276 -3142
rect 30336 -3190 30348 -3142
rect 30264 -3196 30348 -3190
rect 30276 -3230 30336 -3196
rect 30276 -3296 30336 -3290
rect 24944 -3768 25008 -3468
rect 25968 -3640 26160 -3424
rect 25968 -3768 26496 -3640
rect 24944 -3832 26496 -3768
rect 24364 -4236 26156 -4044
rect 24364 -4312 24556 -4236
rect 23624 -4504 24556 -4312
rect 24944 -4412 25008 -4236
rect 25964 -4496 26156 -4236
rect 7904 -7156 8096 -5644
rect 24944 -6412 25008 -4968
rect 25072 -7244 25264 -4608
rect 26304 -5304 26496 -3832
rect 36286 -4496 36346 -4484
rect 30264 -4542 30348 -4536
rect 30264 -4590 30276 -4542
rect 30336 -4590 30348 -4542
rect 30264 -4596 30348 -4590
rect 36286 -4544 36292 -4496
rect 36340 -4544 36346 -4496
rect 30276 -4630 30336 -4596
rect 30276 -4696 30336 -4690
rect 35688 -4892 35864 -4886
rect 35182 -4898 35688 -4892
rect 35182 -5062 35194 -4898
rect 35358 -5062 35688 -4898
rect 35182 -5068 35688 -5062
rect 35688 -5074 35864 -5068
rect 25712 -5496 26496 -5304
rect 31592 -5430 31652 -5418
rect 36286 -5430 36346 -4544
rect 31592 -5490 31598 -5430
rect 31646 -5490 36346 -5430
rect 25712 -5704 25904 -5496
rect 31592 -5502 31652 -5490
rect 30264 -5982 30348 -5976
rect 30264 -6030 30276 -5982
rect 30336 -6030 30348 -5982
rect 30264 -6036 30348 -6030
rect 30276 -6070 30336 -6036
rect 30276 -6136 30336 -6130
rect 24678 -7250 25264 -7244
rect 24678 -7430 24690 -7250
rect 24870 -7430 25264 -7250
rect 24678 -7436 25264 -7430
rect 22888 -8092 23012 -8028
rect 22888 -8412 22952 -8092
rect 25712 -9245 25904 -6444
rect 30264 -7382 30348 -7376
rect 30264 -7430 30276 -7382
rect 30336 -7430 30348 -7382
rect 30264 -7436 30348 -7430
rect 30276 -7470 30336 -7436
rect 30276 -7536 30336 -7530
rect 30264 -8782 30348 -8776
rect 30264 -8830 30276 -8782
rect 30336 -8830 30348 -8782
rect 30264 -8836 30348 -8830
rect 30276 -8870 30336 -8836
rect 30276 -8936 30336 -8930
rect 25712 -9260 29021 -9245
rect 25712 -9376 28576 -9260
rect 25725 -9380 28576 -9376
rect 28796 -9380 29021 -9260
rect 25725 -9395 29021 -9380
rect 29171 -9395 29177 -9245
rect 20892 -15784 21084 -14744
rect 20684 -15976 21084 -15784
<< via1 >>
rect 29856 -1848 30032 -1672
rect 36456 -1868 36632 -1692
rect 30276 -3290 30336 -3230
rect 30276 -4690 30336 -4630
rect 35688 -5068 35864 -4892
rect 30276 -6130 30336 -6070
rect 30276 -7530 30336 -7470
rect 30276 -8930 30336 -8870
rect 29021 -9395 29171 -9245
<< metal2 >>
rect 29856 -1672 30032 -1666
rect 29856 -1957 30032 -1848
rect 36456 -1692 36632 -1686
rect 36456 -1937 36632 -1868
rect 29852 -2123 29861 -1957
rect 30027 -2123 30036 -1957
rect 36452 -2103 36461 -1937
rect 36627 -2103 36636 -1937
rect 36456 -2108 36632 -2103
rect 29856 -2128 30032 -2123
rect 30270 -3290 30276 -3230
rect 30336 -3290 30342 -3230
rect 30276 -3330 30336 -3290
rect 30117 -3390 30126 -3330
rect 30182 -3390 30336 -3330
rect 30270 -4690 30276 -4630
rect 30336 -4690 30342 -4630
rect 30276 -4730 30336 -4690
rect 30117 -4790 30126 -4730
rect 30182 -4790 30336 -4730
rect 35921 -4892 36087 -4888
rect 35682 -5068 35688 -4892
rect 35864 -4897 36092 -4892
rect 35864 -5063 35921 -4897
rect 36087 -5063 36092 -4897
rect 35864 -5068 36092 -5063
rect 35921 -5072 36087 -5068
rect 30270 -6130 30276 -6070
rect 30336 -6130 30342 -6070
rect 30276 -6170 30336 -6130
rect 30117 -6230 30126 -6170
rect 30182 -6230 30336 -6170
rect 30270 -7530 30276 -7470
rect 30336 -7530 30342 -7470
rect 30276 -7570 30336 -7530
rect 30117 -7630 30126 -7570
rect 30182 -7630 30336 -7570
rect 30270 -8930 30276 -8870
rect 30336 -8930 30342 -8870
rect 30276 -8970 30336 -8930
rect 30117 -9030 30126 -8970
rect 30182 -9030 30336 -8970
rect 29021 -9245 29171 -9239
rect 29171 -9395 29351 -9245
rect 29491 -9395 29500 -9245
rect 29021 -9401 29171 -9395
<< via2 >>
rect 29861 -2123 30027 -1957
rect 36461 -2103 36627 -1937
rect 30126 -3390 30182 -3330
rect 30126 -4790 30182 -4730
rect 35921 -5063 36087 -4897
rect 30126 -6230 30182 -6170
rect 30126 -7630 30182 -7570
rect 30126 -9030 30182 -8970
rect 29351 -9395 29491 -9245
<< metal3 >>
rect 36456 -1937 36632 -1932
rect 29856 -1957 30032 -1952
rect 29856 -2123 29861 -1957
rect 30027 -2123 30032 -1957
rect 29316 -9240 29492 -2692
rect 29856 -8652 30032 -2123
rect 36456 -2103 36461 -1937
rect 36627 -2103 36632 -1937
rect 30121 -3330 30187 -3325
rect 30121 -3390 30126 -3330
rect 30182 -3390 31486 -3330
rect 30121 -3395 30187 -3390
rect 30121 -4730 30187 -4725
rect 30121 -4790 30126 -4730
rect 30182 -4790 31506 -4730
rect 30121 -4795 30187 -4790
rect 35916 -4897 36092 -2852
rect 36456 -3888 36632 -2103
rect 35916 -5063 35921 -4897
rect 36087 -5063 36092 -4897
rect 35916 -5068 36092 -5063
rect 30121 -6170 30187 -6165
rect 30121 -6230 30126 -6170
rect 30182 -6230 31606 -6170
rect 30121 -6235 30187 -6230
rect 30121 -7570 30187 -7565
rect 30121 -7630 30126 -7570
rect 30182 -7630 31566 -7570
rect 30121 -7635 30187 -7630
rect 30121 -8970 30187 -8965
rect 30121 -9030 30126 -8970
rect 30182 -9030 31626 -8970
rect 30121 -9035 30187 -9030
rect 29316 -9245 29496 -9240
rect 29316 -9395 29351 -9245
rect 29491 -9395 29583 -9245
rect 29731 -9395 29737 -9245
rect 29316 -9400 29496 -9395
rect 29316 -9408 29492 -9400
<< via3 >>
rect 29583 -9395 29731 -9245
<< metal4 >>
rect 29582 -9245 29732 -9244
rect 31921 -9245 32071 -3695
rect 29582 -9395 29583 -9245
rect 29731 -9395 32071 -9245
rect 29582 -9396 29732 -9395
use JNWTR_CAPX1  JNWTR_CAPX1_0 ../JNW_TR_SKY130A
timestamp 1744633932
transform 0 1 31236 1 0 -9720
box 0 0 1080 1080
use JNWTR_IVX4_CV  JNWTR_IVX4_CV_0 ../JNW_TR_SKY130A
timestamp 1744633932
transform 1 0 28686 0 1 -8680
box -150 -120 2130 920
use JNWTR_IVX4_CV  JNWTR_IVX4_CV_1
timestamp 1744633932
transform 1 0 28686 0 1 -4380
box -150 -120 2130 920
use JNWTR_IVX4_CV  JNWTR_IVX4_CV_2
timestamp 1744633932
transform 1 0 28686 0 1 -7180
box -150 -120 2130 920
use JNWTR_IVX4_CV  JNWTR_IVX4_CV_3
timestamp 1744633932
transform 1 0 28686 0 1 -5880
box -150 -120 2130 920
use JNWTR_IVX4_CV  JNWTR_IVX4_CV_4
timestamp 1744633932
transform 1 0 28686 0 1 -2980
box -150 -120 2130 920
use JNW_VIS_TI  x2 ../JNW_GR02_SKY130A
timestamp 1745488532
transform 1 0 14388 0 1 1400
box -9344 -19400 9900 -2398
use JNWTR_CAPX1  x7
timestamp 1744633932
transform 0 -1 32316 1 0 -3800
box 0 0 1080 1080
use JNWATR_NCH_8C1F2  x8 ../JNW_ATR_SKY130A
timestamp 1744633932
transform 1 0 24784 0 1 -7072
box -184 -128 1592 928
use JNWATR_NCH_12C1F2  x9 ../JNW_ATR_SKY130A
timestamp 1744633932
transform 1 0 24784 0 1 -5072
box -184 -128 1848 928
use JNWTR_IVX4_CV  x10
timestamp 1744633932
transform 1 0 35286 0 1 -3080
box -150 -120 2130 920
use JNWATR_NCH_8C1F2  x11
timestamp 1744633932
transform 1 0 24784 0 1 -6272
box -184 -128 1592 928
use JNWATR_PCH_12C1F2  x12 ../JNW_ATR_SKY130A
timestamp 1744633932
transform 1 0 24784 0 1 -3672
box -184 -128 1848 928
use JNWATR_PCH_12C1F2  x13
timestamp 1744633932
transform 1 0 24784 0 1 -2872
box -184 -128 1848 928
use JNWTR_IVX4_CV  x14
timestamp 1744633932
transform 1 0 35286 0 1 -4420
box -150 -120 2130 920
use JNWTR_CAPX1  x15
timestamp 1744633932
transform 0 -1 32316 1 0 -5300
box 0 0 1080 1080
use JNWTR_CAPX1  x16
timestamp 1744633932
transform 0 -1 32316 1 0 -6800
box 0 0 1080 1080
use JNWTR_CAPX1  x17
timestamp 1744633932
transform 0 -1 32316 1 0 -8300
box 0 0 1080 1080
<< labels >>
flabel locali 24688 -10216 26686 -10024 0 FreeSans 1600 0 0 0 VSS
port 0 nsew
flabel metal1 22948 -8092 23012 -8028 0 FreeSans 1600 0 0 0 PWR_UP
port 2 nsew
flabel locali 29060 -1196 29252 -1004 0 FreeSans 1600 0 0 0 VDD
port 3 nsew
flabel locali 36006 -2010 36066 -1950 0 FreeSans 1600 0 0 0 VOUT
port 1 nsew
flabel metal1 7904 -5836 8096 -5644 0 FreeSans 1600 0 0 0 VREF
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 34124 12080
<< end >>
