magic
tech sky130A
magscale 1 2
timestamp 1744473896
<< checkpaint >>
rect -6764 12310 -4243 14709
rect -16108 11793 5656 12310
rect 8389 11793 10910 13786
rect -16108 -7212 20890 11793
rect -6387 -13325 20890 -7212
rect -6387 -16983 5528 -13325
rect -6387 -17807 -3866 -16983
<< locali >>
rect 15616 4416 17408 4544
rect 14840 4066 14900 4258
rect 15616 4160 15680 4416
rect 17344 4096 17408 4416
rect 18082 4170 18142 4386
rect 14840 4064 14848 4066
<< viali >>
rect 14840 4258 14900 4318
rect 18082 4386 18142 4446
<< metal1 >>
rect -14100 4892 -1456 5084
rect 988 3636 2854 3700
rect 3732 3232 3924 5744
rect 19264 4800 19392 6720
rect 14807 4673 19392 4800
rect 14807 4318 14934 4673
rect 14976 4672 19392 4673
rect 18076 4452 18148 4458
rect 18070 4392 18076 4452
rect 18148 4392 18154 4452
rect 18070 4386 18082 4392
rect 18142 4386 18154 4392
rect 18070 4380 18154 4386
rect 14807 4289 14840 4318
rect 14828 4258 14840 4289
rect 14900 4289 14934 4318
rect 14900 4258 14912 4289
rect 14828 4252 14912 4258
rect 10817 3455 10944 3461
rect 10944 3328 11647 3455
rect 10817 3322 10944 3328
rect 3732 3040 12000 3232
rect 10817 2944 10944 2950
rect 3777 2942 10817 2943
rect 2307 2819 10817 2942
rect 2307 -6850 2430 2819
rect 3777 2817 10817 2819
rect 10817 2811 10944 2817
rect -5117 -6973 2430 -6850
rect -5117 -6979 -4994 -6973
rect -5117 -7108 -4994 -7102
<< via1 >>
rect 18076 4446 18148 4452
rect 18076 4392 18082 4446
rect 18082 4392 18142 4446
rect 18142 4392 18148 4446
rect 10817 3328 10944 3455
rect 10817 2817 10944 2944
rect -5117 -7102 -4994 -6979
<< metal2 >>
rect 13441 4865 18176 4992
rect 10811 3328 10817 3455
rect 10944 3328 10950 3455
rect 10817 2944 10944 3328
rect 13441 2944 13568 4865
rect 18082 4452 18142 4865
rect 18070 4392 18076 4452
rect 18148 4392 18154 4452
rect 10811 2817 10817 2944
rect 10944 2817 13568 2944
rect -5123 -7102 -5117 -6979
rect -4994 -7102 -4988 -6979
rect -5117 -7234 -4994 -7102
rect -5117 -7366 -4994 -7357
<< via2 >>
rect -5117 -7357 -4994 -7234
<< metal3 >>
rect 15872 4480 18520 4608
rect 15872 3968 16000 4480
rect 15360 3136 15488 3520
rect 17804 3136 17980 4024
rect 18344 3704 18520 4480
rect 15360 3008 17984 3136
rect -5122 -7234 -4989 -7229
rect -5122 -7357 -5117 -7234
rect -4994 -7357 -4989 -7234
rect -5122 -7362 -4989 -7357
rect -5116 -8061 -4993 -7362
use JNW_VIS_ITIME  x1 ../JNW_GR02_SKY130A
timestamp 1744462317
transform 1 0 9649 0 1 12525
box -4352 -24590 9981 -1992
use JNW_VIS_TI  x2 ../JNW_GR02_SKY130A
timestamp 1744467493
transform 1 0 -5504 0 1 13448
box -9344 -19400 9900 -2398
use JNWTR_DFTSPCX1_CV  x3 ../JNW_TR_SKY130A
timestamp 1744464884
transform 1 0 14690 0 1 3314
box -150 -120 2130 1080
use JNWTR_DFTSPCX1_CV  x4
timestamp 1744464884
transform 1 0 17174 0 1 3320
box -150 -120 2130 1080
use dig  x5 ../JNW_GR02_SKY130A
timestamp 1744314437
transform 1 0 -5127 0 1 -16547
box 0 824 9395 10464
<< properties >>
string FIXED_BBOX 0 0 22267 11539
<< end >>
