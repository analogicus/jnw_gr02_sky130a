** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_GR02_SKY130A/TB_JNW_VIS_TI.sch
**.subckt TB_JNW_VIS_TI VDD VSS VREF I_TEMP PWR_UP LPI LPO
*.ipin VDD
*.ipin VSS
*.opin VREF
*.opin I_TEMP
*.ipin PWR_UP
*.opin LPI
*.opin LPO
x1 I_TEMP VDD VREF LPO LPI PWR_UP VSS JNW_VIS_TI
**** begin user architecture code



.param mc_mm_switch=0
.param mc_pr_switch=0
.include tt.spi
*.include ss.spi
.option gmin=1e-15
.lib ../../../tech/ngspice/temperature.spi Tl
.lib ../../../tech/ngspice/supply.spi Vl
.include ../../../../cpdk/ngspice/ideal_circuits.spi
.include /home/domen/pro/aicex/ip/cpdk/ngspice/tian_subckt.lib

X999 LPI LPO loopgainprobe

VSS  VSS  0     dc 0
VDD  VDD VSS dc 1.8
VPUP PWR_UP VSS PULSE ( 0 1.8 10NS 1PS 1PS 10NS 1S 1)
VSENS I_TEMP VSS dc 0.6


.option temp = 27
.option savecurrents
.save all
.control

.IC V(LPO)=0.5
optran 0 0 0 10n 100u 0
op
write TB_JNW_VIS_TI.raw
exit
.endc
.end



**** end user architecture code
**.ends

* expanding   symbol:  JNW_GR02_SKY130A/JNW_VIS_TI.sym # of pins=7
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_GR02_SKY130A/JNW_VIS_TI.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_GR02_SKY130A/JNW_VIS_TI.sch
.subckt JNW_VIS_TI I_TEMP VDD VREF LPO LPI PWR_UP VSS
*.ipin VSS
*.opin VREF
*.ipin PWR_UP
*.opin LPI
*.opin LPO
*.ipin VDD
*.opin I_TEMP
XQ1<0> VSS VSS VIN sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1 mult=1
XQ2<0> VSS VSS VD2 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=8 mult=8
x7 VDD VIN VIP VSS LPO JNW_VIS_OTA
x11<0> LPI PWR_UP VSS VSS JNWATR_NCH_4C5F0
x11<1> LPI PWR_UP VSS VSS JNWATR_NCH_4C5F0
x1<0> LPI VSS JNWTR_CAPX1
x1<1> LPI VSS JNWTR_CAPX1
x1<2> LPI VSS JNWTR_CAPX1
x1<3> LPI VSS JNWTR_CAPX1
x1<4> LPI VSS JNWTR_CAPX1
x1<5> LPI VSS JNWTR_CAPX1
x1<6> LPI VSS JNWTR_CAPX1
x1<7> LPI VSS JNWTR_CAPX1
x1<8> LPI VSS JNWTR_CAPX1
x1<9> LPI VSS JNWTR_CAPX1
x1<10> LPI VSS JNWTR_CAPX1
x1<11> LPI VSS JNWTR_CAPX1
x1<12> LPI VSS JNWTR_CAPX1
x1<13> LPI VSS JNWTR_CAPX1
x1<14> LPI VSS JNWTR_CAPX1
x1<15> LPI VSS JNWTR_CAPX1
x1<16> LPI VSS JNWTR_CAPX1
x1<17> LPI VSS JNWTR_CAPX1
x1<18> LPI VSS JNWTR_CAPX1
x1<19> LPI VSS JNWTR_CAPX1
x9 V_MEAS1 LPI VSS VSS JNWATR_NCH_12C5F0
x2<0> V_MEAS2 V_MEAS1 VDD VDD JNWATR_PCH_4C5F0
x2<1> V_MEAS2 V_MEAS1 VDD VDD JNWATR_PCH_4C5F0
x2<2> V_MEAS2 V_MEAS1 VDD VDD JNWATR_PCH_4C5F0
x3<0> V_MEAS1 V_MEAS3 V_MEAS2 V_MEAS2 JNWATR_PCH_4C5F0
x3<1> V_MEAS1 V_MEAS3 V_MEAS2 V_MEAS2 JNWATR_PCH_4C5F0
x3<2> V_MEAS1 V_MEAS3 V_MEAS2 V_MEAS2 JNWATR_PCH_4C5F0
x4<0> V_MEAS4 V_MEAS1 VDD VDD JNWATR_PCH_4C5F0
x4<1> V_MEAS4 V_MEAS1 VDD VDD JNWATR_PCH_4C5F0
x4<2> V_MEAS4 V_MEAS1 VDD VDD JNWATR_PCH_4C5F0
x5<0> VREF V_MEAS3 V_MEAS4 V_MEAS4 JNWATR_PCH_4C5F0
x5<1> VREF V_MEAS3 V_MEAS4 V_MEAS4 JNWATR_PCH_4C5F0
x5<2> VREF V_MEAS3 V_MEAS4 V_MEAS4 JNWATR_PCH_4C5F0
x15 V_MEAS3 V_MEAS3 VDD VDD JNWATR_PCH_2C5F0
x6<0> net2<2> V_MEAS1 VDD VDD JNWATR_PCH_4C5F0
x6<1> net2<1> V_MEAS1 VDD VDD JNWATR_PCH_4C5F0
x6<2> net2<0> V_MEAS1 VDD VDD JNWATR_PCH_4C5F0
x8<0> VSS V_MEAS3 net2<2> net2<2> JNWATR_PCH_4C5F0
x8<1> VSS V_MEAS3 net2<1> net2<1> JNWATR_PCH_4C5F0
x8<2> VSS V_MEAS3 net2<0> net2<0> JNWATR_PCH_4C5F0
x7<0> net1<2> V_MEAS1 VDD VDD JNWATR_PCH_4C5F0
x7<1> net1<1> V_MEAS1 VDD VDD JNWATR_PCH_4C5F0
x7<2> net1<0> V_MEAS1 VDD VDD JNWATR_PCH_4C5F0
x10<0> VIN V_MEAS3 net1<2> net1<2> JNWATR_PCH_4C5F0
x10<1> VIN V_MEAS3 net1<1> net1<1> JNWATR_PCH_4C5F0
x10<2> VIN V_MEAS3 net1<0> net1<0> JNWATR_PCH_4C5F0
x14 net3 VREF VSS JNWTR_RPPO2
x12<0> net6<1> net3 VSS JNWTR_RPPO2
x12<1> net6<0> net3 VSS JNWTR_RPPO2
x13<0> VD2 VIP VSS JNWTR_RPPO2
x13<1> VD2 VIP VSS JNWTR_RPPO2
x13<2> VD2 VIP VSS JNWTR_RPPO2
x13<3> VD2 VIP VSS JNWTR_RPPO2
x9<0> net4<1> V_MEAS3 VSS JNWTR_RPPO2
x9<1> net4<0> V_MEAS3 VSS JNWTR_RPPO2
x15<0> VSS net4<1> VSS JNWTR_RPPO2
x15<1> VSS net4<0> VSS JNWTR_RPPO2
x2 net5 V_MEAS1 VDD VDD JNWATR_PCH_2C5F0
x14<0> VIP net6<1> VSS JNWTR_RPPO2
x14<1> VIP net6<0> VSS JNWTR_RPPO2
x16<0> I_TEMP V_MEAS3 net5 net5 JNWATR_PCH_4C5F0
x16<1> I_TEMP V_MEAS3 net5 net5 JNWATR_PCH_4C5F0
x16<2> I_TEMP V_MEAS3 net5 net5 JNWATR_PCH_4C5F0
.ends


* expanding   symbol:  JNW_GR02_SKY130A/JNW_VIS_OTA.sym # of pins=5
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_GR02_SKY130A/JNW_VIS_OTA.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_GR02_SKY130A/JNW_VIS_OTA.sch
.subckt JNW_VIS_OTA VDD VIN VIP VSS VOUT
*.ipin VDD
*.ipin VIP
*.ipin VIN
*.ipin VSS
*.opin VOUT
x7<0> V2 VIP VOP VDD JNWATR_PCH_12C1F2
x7<1> V2 VIP VOP VDD JNWATR_PCH_12C1F2
x7<2> V2 VIP VOP VDD JNWATR_PCH_12C1F2
x7<3> V2 VIP VOP VDD JNWATR_PCH_12C1F2
x1<0> V1 VIN VOP VDD JNWATR_PCH_12C1F2
x1<1> V1 VIN VOP VDD JNWATR_PCH_12C1F2
x1<2> V1 VIN VOP VDD JNWATR_PCH_12C1F2
x1<3> V1 VIN VOP VDD JNWATR_PCH_12C1F2
x10 VOUT V1 VSS VSS JNWATR_NCH_12C5F0
x5 V2 V2 VSS VSS JNWATR_NCH_12C5F0
x2 net1 V2 VSS VSS JNWATR_NCH_12C5F0
x3 V1 V1 VSS VSS JNWATR_NCH_12C5F0
x2<0> VOUT net1 VDD VDD JNWATR_PCH_12C5F0
x2<1> VOUT net1 VDD VDD JNWATR_PCH_12C5F0
x2<2> VOUT net1 VDD VDD JNWATR_PCH_12C5F0
x2<3> VOUT net1 VDD VDD JNWATR_PCH_12C5F0
x3<0> net1 net1 VDD VDD JNWATR_PCH_12C5F0
x3<1> net1 net1 VDD VDD JNWATR_PCH_12C5F0
x3<2> net1 net1 VDD VDD JNWATR_PCH_12C5F0
x3<3> net1 net1 VDD VDD JNWATR_PCH_12C5F0
x6 net3 net2 VSS JNWTR_RPPO2
x8<0> VSS net3 VSS JNWTR_RPPO2
x8<1> VSS net3 VSS JNWTR_RPPO2
x13 net2 net2 VDD VDD JNWATR_PCH_12C5F0
x14 VOP net2 VDD VDD JNWATR_PCH_12C5F0
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sch
.subckt JNWATR_NCH_4C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.94 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_CAPX1.sym # of pins=2
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sch
.subckt JNWTR_CAPX1 A B
*.iopin A
*.iopin B
XC1 B A sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_12C5F0.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_12C5F0.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_12C5F0.sch
.subckt JNWATR_NCH_12C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.94 W=8.32 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sch
.subckt JNWATR_PCH_4C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.94 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_2C5F0.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_2C5F0.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_2C5F0.sch
.subckt JNWATR_PCH_2C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.94 W=1.92 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RPPO2.sym # of pins=3
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO2.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO2.sch
.subckt JNWTR_RPPO2 N P B
*.iopin P
*.iopin N
*.iopin B
XXA1 N P B JNWTR_RES2
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_12C1F2.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_12C1F2.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_12C1F2.sch
.subckt JNWATR_PCH_12C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.22 W=8.32 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_12C5F0.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_12C5F0.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_12C5F0.sch
.subckt JNWATR_PCH_12C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.94 W=8.32 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RES2.sym # of pins=3
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RES2.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RES2.sch
.subckt JNWTR_RES2 N P B
*.iopin N
*.iopin P
*.iopin B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_1 P INT_0 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
.ends

.end
