magic
tech sky130A
magscale 1 2
timestamp 1744314437
<< viali >>
rect 2881 9129 2915 9163
rect 7665 9129 7699 9163
rect 3893 8993 3927 9027
rect 4629 8993 4663 9027
rect 4721 8993 4755 9027
rect 4905 8993 4939 9027
rect 7205 8993 7239 9027
rect 1409 8925 1443 8959
rect 3065 8925 3099 8959
rect 3157 8925 3191 8959
rect 3525 8925 3559 8959
rect 3617 8925 3651 8959
rect 4077 8925 4111 8959
rect 4169 8925 4203 8959
rect 4445 8925 4479 8959
rect 5549 8925 5583 8959
rect 7021 8925 7055 8959
rect 7481 8925 7515 8959
rect 5457 8857 5491 8891
rect 7113 8857 7147 8891
rect 1593 8789 1627 8823
rect 3433 8789 3467 8823
rect 3893 8789 3927 8823
rect 4261 8789 4295 8823
rect 6193 8789 6227 8823
rect 6653 8789 6687 8823
rect 4077 8585 4111 8619
rect 6745 8585 6779 8619
rect 4353 8517 4387 8551
rect 6837 8517 6871 8551
rect 2513 8449 2547 8483
rect 2697 8449 2731 8483
rect 2973 8449 3007 8483
rect 3709 8449 3743 8483
rect 3801 8449 3835 8483
rect 3985 8449 4019 8483
rect 4261 8449 4295 8483
rect 4445 8449 4479 8483
rect 4629 8449 4663 8483
rect 4813 8449 4847 8483
rect 5457 8449 5491 8483
rect 5641 8449 5675 8483
rect 6561 8381 6595 8415
rect 7297 8381 7331 8415
rect 2697 8313 2731 8347
rect 3985 8313 4019 8347
rect 7205 8313 7239 8347
rect 3433 8245 3467 8279
rect 6193 8245 6227 8279
rect 7941 8245 7975 8279
rect 3985 8041 4019 8075
rect 6561 8041 6595 8075
rect 2973 7973 3007 8007
rect 3525 7905 3559 7939
rect 4629 7905 4663 7939
rect 1593 7837 1627 7871
rect 3157 7837 3191 7871
rect 3617 7837 3651 7871
rect 6469 7837 6503 7871
rect 7941 7837 7975 7871
rect 1860 7769 1894 7803
rect 4721 7769 4755 7803
rect 7674 7769 7708 7803
rect 5365 7497 5399 7531
rect 7757 7497 7791 7531
rect 4252 7429 4286 7463
rect 6622 7429 6656 7463
rect 2513 7361 2547 7395
rect 2780 7361 2814 7395
rect 5825 7361 5859 7395
rect 6377 7361 6411 7395
rect 3985 7293 4019 7327
rect 5641 7293 5675 7327
rect 5733 7293 5767 7327
rect 3893 7157 3927 7191
rect 6193 7157 6227 7191
rect 5273 6953 5307 6987
rect 2145 6817 2179 6851
rect 5457 6817 5491 6851
rect 7757 6817 7791 6851
rect 1869 6749 1903 6783
rect 1961 6749 1995 6783
rect 2329 6749 2363 6783
rect 2973 6749 3007 6783
rect 3617 6749 3651 6783
rect 3893 6749 3927 6783
rect 5365 6749 5399 6783
rect 5549 6749 5583 6783
rect 5733 6749 5767 6783
rect 2881 6681 2915 6715
rect 4138 6681 4172 6715
rect 6000 6681 6034 6715
rect 2145 6613 2179 6647
rect 7113 6613 7147 6647
rect 7205 6613 7239 6647
rect 7573 6613 7607 6647
rect 7665 6613 7699 6647
rect 2605 6409 2639 6443
rect 4261 6409 4295 6443
rect 4429 6409 4463 6443
rect 6193 6409 6227 6443
rect 2421 6341 2455 6375
rect 4629 6341 4663 6375
rect 2697 6273 2731 6307
rect 3056 6273 3090 6307
rect 5181 6273 5215 6307
rect 6377 6273 6411 6307
rect 6644 6273 6678 6307
rect 2789 6205 2823 6239
rect 5089 6205 5123 6239
rect 5273 6205 5307 6239
rect 5365 6205 5399 6239
rect 5641 6205 5675 6239
rect 2421 6137 2455 6171
rect 4169 6137 4203 6171
rect 4445 6069 4479 6103
rect 4905 6069 4939 6103
rect 7757 6069 7791 6103
rect 5365 5865 5399 5899
rect 6101 5865 6135 5899
rect 6837 5865 6871 5899
rect 7849 5865 7883 5899
rect 3617 5797 3651 5831
rect 6653 5729 6687 5763
rect 7389 5729 7423 5763
rect 3157 5661 3191 5695
rect 3433 5661 3467 5695
rect 7665 5661 7699 5695
rect 3249 5593 3283 5627
rect 4077 5593 4111 5627
rect 4813 5321 4847 5355
rect 4997 5321 5031 5355
rect 6745 5321 6779 5355
rect 7205 5321 7239 5355
rect 2697 5253 2731 5287
rect 2913 5253 2947 5287
rect 5181 5253 5215 5287
rect 3341 5185 3375 5219
rect 5089 5185 5123 5219
rect 6837 5185 6871 5219
rect 7757 5185 7791 5219
rect 3617 5117 3651 5151
rect 4077 5117 4111 5151
rect 5641 5117 5675 5151
rect 7021 5117 7055 5151
rect 3065 5049 3099 5083
rect 5365 5049 5399 5083
rect 6377 5049 6411 5083
rect 2881 4981 2915 5015
rect 3157 4981 3191 5015
rect 3525 4981 3559 5015
rect 4629 4981 4663 5015
rect 6193 4981 6227 5015
rect 3617 4777 3651 4811
rect 5549 4777 5583 4811
rect 7481 4777 7515 4811
rect 7849 4777 7883 4811
rect 2605 4709 2639 4743
rect 2881 4641 2915 4675
rect 4169 4641 4203 4675
rect 3065 4573 3099 4607
rect 3801 4573 3835 4607
rect 4425 4573 4459 4607
rect 5733 4573 5767 4607
rect 6101 4573 6135 4607
rect 6357 4573 6391 4607
rect 7665 4573 7699 4607
rect 3893 4505 3927 4539
rect 4077 4505 4111 4539
rect 2421 4437 2455 4471
rect 3801 4437 3835 4471
rect 5917 4437 5951 4471
rect 3801 4233 3835 4267
rect 4445 4165 4479 4199
rect 2688 4097 2722 4131
rect 4353 4097 4387 4131
rect 6633 4097 6667 4131
rect 2421 4029 2455 4063
rect 4261 4029 4295 4063
rect 6377 4029 6411 4063
rect 5733 3893 5767 3927
rect 7757 3893 7791 3927
rect 5273 3689 5307 3723
rect 7389 3689 7423 3723
rect 7849 3689 7883 3723
rect 3617 3621 3651 3655
rect 2237 3553 2271 3587
rect 3893 3553 3927 3587
rect 2504 3485 2538 3519
rect 5457 3485 5491 3519
rect 6009 3485 6043 3519
rect 7665 3485 7699 3519
rect 4138 3417 4172 3451
rect 6254 3417 6288 3451
rect 2973 3145 3007 3179
rect 5365 3145 5399 3179
rect 7757 3145 7791 3179
rect 4629 3077 4663 3111
rect 5917 3077 5951 3111
rect 3065 3009 3099 3043
rect 3157 3009 3191 3043
rect 3341 3009 3375 3043
rect 5825 3009 5859 3043
rect 6377 3009 6411 3043
rect 6644 3009 6678 3043
rect 2697 2941 2731 2975
rect 4077 2941 4111 2975
rect 4813 2941 4847 2975
rect 6009 2941 6043 2975
rect 5457 2873 5491 2907
rect 3893 2805 3927 2839
rect 3433 2601 3467 2635
rect 3893 2601 3927 2635
rect 5917 2601 5951 2635
rect 6653 2601 6687 2635
rect 7849 2601 7883 2635
rect 3617 2533 3651 2567
rect 5365 2465 5399 2499
rect 7113 2465 7147 2499
rect 7205 2465 7239 2499
rect 3157 2397 3191 2431
rect 4077 2397 4111 2431
rect 4353 2397 4387 2431
rect 4537 2397 4571 2431
rect 7665 2397 7699 2431
rect 3249 2329 3283 2363
rect 3465 2329 3499 2363
rect 7021 2329 7055 2363
rect 2973 2261 3007 2295
rect 4261 2261 4295 2295
rect 5089 2261 5123 2295
rect 5457 2261 5491 2295
rect 5549 2261 5583 2295
<< metal1 >>
rect 3050 9324 3056 9376
rect 3108 9364 3114 9376
rect 5534 9364 5540 9376
rect 3108 9336 5540 9364
rect 3108 9324 3114 9336
rect 5534 9324 5540 9336
rect 5592 9324 5598 9376
rect 1104 9274 8280 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 8280 9274
rect 1104 9200 8280 9222
rect 2869 9163 2927 9169
rect 2869 9129 2881 9163
rect 2915 9160 2927 9163
rect 6914 9160 6920 9172
rect 2915 9132 6920 9160
rect 2915 9129 2927 9132
rect 2869 9123 2927 9129
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 7650 9120 7656 9172
rect 7708 9120 7714 9172
rect 3528 9064 4752 9092
rect 842 8916 848 8968
rect 900 8956 906 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 900 8928 1409 8956
rect 900 8916 906 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 3050 8916 3056 8968
rect 3108 8916 3114 8968
rect 3145 8959 3203 8965
rect 3145 8925 3157 8959
rect 3191 8956 3203 8959
rect 3418 8956 3424 8968
rect 3191 8928 3424 8956
rect 3191 8925 3203 8928
rect 3145 8919 3203 8925
rect 3418 8916 3424 8928
rect 3476 8916 3482 8968
rect 3528 8965 3556 9064
rect 3694 8984 3700 9036
rect 3752 9024 3758 9036
rect 4724 9033 4752 9064
rect 4908 9064 7512 9092
rect 4908 9033 4936 9064
rect 3881 9027 3939 9033
rect 3881 9024 3893 9027
rect 3752 8996 3893 9024
rect 3752 8984 3758 8996
rect 3881 8993 3893 8996
rect 3927 8993 3939 9027
rect 4617 9027 4675 9033
rect 4617 9024 4629 9027
rect 3881 8987 3939 8993
rect 3988 8996 4629 9024
rect 3513 8959 3571 8965
rect 3513 8925 3525 8959
rect 3559 8925 3571 8959
rect 3513 8919 3571 8925
rect 3605 8959 3663 8965
rect 3605 8925 3617 8959
rect 3651 8956 3663 8959
rect 3786 8956 3792 8968
rect 3651 8928 3792 8956
rect 3651 8925 3663 8928
rect 3605 8919 3663 8925
rect 3786 8916 3792 8928
rect 3844 8956 3850 8968
rect 3988 8956 4016 8996
rect 4617 8993 4629 8996
rect 4663 8993 4675 9027
rect 4617 8987 4675 8993
rect 4709 9027 4767 9033
rect 4709 8993 4721 9027
rect 4755 9024 4767 9027
rect 4893 9027 4951 9033
rect 4755 8996 4844 9024
rect 4755 8993 4767 8996
rect 4709 8987 4767 8993
rect 3844 8928 4016 8956
rect 3844 8916 3850 8928
rect 4062 8916 4068 8968
rect 4120 8916 4126 8968
rect 4154 8916 4160 8968
rect 4212 8916 4218 8968
rect 4433 8959 4491 8965
rect 4433 8925 4445 8959
rect 4479 8925 4491 8959
rect 4816 8956 4844 8996
rect 4893 8993 4905 9027
rect 4939 8993 4951 9027
rect 4893 8987 4951 8993
rect 5442 8984 5448 9036
rect 5500 9024 5506 9036
rect 5500 8996 7052 9024
rect 5500 8984 5506 8996
rect 5258 8956 5264 8968
rect 4816 8928 5264 8956
rect 4433 8919 4491 8925
rect 2958 8888 2964 8900
rect 2746 8860 2964 8888
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 2746 8820 2774 8860
rect 2958 8848 2964 8860
rect 3016 8848 3022 8900
rect 4448 8888 4476 8919
rect 5258 8916 5264 8928
rect 5316 8916 5322 8968
rect 5534 8916 5540 8968
rect 5592 8916 5598 8968
rect 7024 8965 7052 8996
rect 7098 8984 7104 9036
rect 7156 9024 7162 9036
rect 7193 9027 7251 9033
rect 7193 9024 7205 9027
rect 7156 8996 7205 9024
rect 7156 8984 7162 8996
rect 7193 8993 7205 8996
rect 7239 8993 7251 9027
rect 7193 8987 7251 8993
rect 7484 8968 7512 9064
rect 7009 8959 7067 8965
rect 7009 8925 7021 8959
rect 7055 8925 7067 8959
rect 7009 8919 7067 8925
rect 7466 8916 7472 8968
rect 7524 8916 7530 8968
rect 3436 8860 4476 8888
rect 5445 8891 5503 8897
rect 3436 8829 3464 8860
rect 5445 8857 5457 8891
rect 5491 8888 5503 8891
rect 7101 8891 7159 8897
rect 7101 8888 7113 8891
rect 5491 8860 7113 8888
rect 5491 8857 5503 8860
rect 5445 8851 5503 8857
rect 7101 8857 7113 8860
rect 7147 8857 7159 8891
rect 7101 8851 7159 8857
rect 1627 8792 2774 8820
rect 3421 8823 3479 8829
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 3421 8789 3433 8823
rect 3467 8789 3479 8823
rect 3421 8783 3479 8789
rect 3881 8823 3939 8829
rect 3881 8789 3893 8823
rect 3927 8820 3939 8823
rect 3970 8820 3976 8832
rect 3927 8792 3976 8820
rect 3927 8789 3939 8792
rect 3881 8783 3939 8789
rect 3970 8780 3976 8792
rect 4028 8780 4034 8832
rect 4249 8823 4307 8829
rect 4249 8789 4261 8823
rect 4295 8820 4307 8823
rect 4614 8820 4620 8832
rect 4295 8792 4620 8820
rect 4295 8789 4307 8792
rect 4249 8783 4307 8789
rect 4614 8780 4620 8792
rect 4672 8780 4678 8832
rect 6178 8780 6184 8832
rect 6236 8780 6242 8832
rect 6638 8780 6644 8832
rect 6696 8780 6702 8832
rect 1104 8730 8280 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 8280 8730
rect 1104 8656 8280 8678
rect 3694 8616 3700 8628
rect 2746 8588 3700 8616
rect 2746 8548 2774 8588
rect 3694 8576 3700 8588
rect 3752 8576 3758 8628
rect 3786 8576 3792 8628
rect 3844 8616 3850 8628
rect 4065 8619 4123 8625
rect 4065 8616 4077 8619
rect 3844 8588 4077 8616
rect 3844 8576 3850 8588
rect 4065 8585 4077 8588
rect 4111 8585 4123 8619
rect 4065 8579 4123 8585
rect 5276 8588 5488 8616
rect 2516 8520 2774 8548
rect 2516 8489 2544 8520
rect 2501 8483 2559 8489
rect 2501 8449 2513 8483
rect 2547 8449 2559 8483
rect 2501 8443 2559 8449
rect 2682 8440 2688 8492
rect 2740 8440 2746 8492
rect 2958 8440 2964 8492
rect 3016 8440 3022 8492
rect 3602 8440 3608 8492
rect 3660 8480 3666 8492
rect 3804 8489 3832 8576
rect 4341 8551 4399 8557
rect 4341 8517 4353 8551
rect 4387 8548 4399 8551
rect 4890 8548 4896 8560
rect 4387 8520 4896 8548
rect 4387 8517 4399 8520
rect 4341 8511 4399 8517
rect 4890 8508 4896 8520
rect 4948 8548 4954 8560
rect 5276 8548 5304 8588
rect 4948 8520 5304 8548
rect 5460 8548 5488 8588
rect 6178 8576 6184 8628
rect 6236 8616 6242 8628
rect 6733 8619 6791 8625
rect 6733 8616 6745 8619
rect 6236 8588 6745 8616
rect 6236 8576 6242 8588
rect 6733 8585 6745 8588
rect 6779 8585 6791 8619
rect 6733 8579 6791 8585
rect 6825 8551 6883 8557
rect 6825 8548 6837 8551
rect 5460 8520 6837 8548
rect 4948 8508 4954 8520
rect 6825 8517 6837 8520
rect 6871 8517 6883 8551
rect 6825 8511 6883 8517
rect 3697 8483 3755 8489
rect 3697 8480 3709 8483
rect 3660 8452 3709 8480
rect 3660 8440 3666 8452
rect 3697 8449 3709 8452
rect 3743 8449 3755 8483
rect 3697 8443 3755 8449
rect 3789 8483 3847 8489
rect 3789 8449 3801 8483
rect 3835 8449 3847 8483
rect 3789 8443 3847 8449
rect 3970 8440 3976 8492
rect 4028 8440 4034 8492
rect 4246 8440 4252 8492
rect 4304 8440 4310 8492
rect 4430 8440 4436 8492
rect 4488 8440 4494 8492
rect 4617 8483 4675 8489
rect 4617 8449 4629 8483
rect 4663 8480 4675 8483
rect 4706 8480 4712 8492
rect 4663 8452 4712 8480
rect 4663 8449 4675 8452
rect 4617 8443 4675 8449
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8480 4859 8483
rect 5258 8480 5264 8492
rect 4847 8452 5264 8480
rect 4847 8449 4859 8452
rect 4801 8443 4859 8449
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 5442 8440 5448 8492
rect 5500 8440 5506 8492
rect 5629 8483 5687 8489
rect 5629 8449 5641 8483
rect 5675 8480 5687 8483
rect 6638 8480 6644 8492
rect 5675 8452 6644 8480
rect 5675 8449 5687 8452
rect 5629 8443 5687 8449
rect 6638 8440 6644 8452
rect 6696 8440 6702 8492
rect 6549 8415 6607 8421
rect 6549 8412 6561 8415
rect 5644 8384 6561 8412
rect 2685 8347 2743 8353
rect 2685 8313 2697 8347
rect 2731 8344 2743 8347
rect 2774 8344 2780 8356
rect 2731 8316 2780 8344
rect 2731 8313 2743 8316
rect 2685 8307 2743 8313
rect 2774 8304 2780 8316
rect 2832 8304 2838 8356
rect 3694 8304 3700 8356
rect 3752 8344 3758 8356
rect 3973 8347 4031 8353
rect 3973 8344 3985 8347
rect 3752 8316 3985 8344
rect 3752 8304 3758 8316
rect 3973 8313 3985 8316
rect 4019 8313 4031 8347
rect 3973 8307 4031 8313
rect 4246 8304 4252 8356
rect 4304 8344 4310 8356
rect 5350 8344 5356 8356
rect 4304 8316 5356 8344
rect 4304 8304 4310 8316
rect 5350 8304 5356 8316
rect 5408 8304 5414 8356
rect 5644 8288 5672 8384
rect 6549 8381 6561 8384
rect 6595 8412 6607 8415
rect 7098 8412 7104 8424
rect 6595 8384 7104 8412
rect 6595 8381 6607 8384
rect 6549 8375 6607 8381
rect 7098 8372 7104 8384
rect 7156 8372 7162 8424
rect 7285 8415 7343 8421
rect 7285 8381 7297 8415
rect 7331 8381 7343 8415
rect 7285 8375 7343 8381
rect 7193 8347 7251 8353
rect 7193 8313 7205 8347
rect 7239 8344 7251 8347
rect 7300 8344 7328 8375
rect 7239 8316 7328 8344
rect 7239 8313 7251 8316
rect 7193 8307 7251 8313
rect 3421 8279 3479 8285
rect 3421 8245 3433 8279
rect 3467 8276 3479 8279
rect 5626 8276 5632 8288
rect 3467 8248 5632 8276
rect 3467 8245 3479 8248
rect 3421 8239 3479 8245
rect 5626 8236 5632 8248
rect 5684 8236 5690 8288
rect 6178 8236 6184 8288
rect 6236 8236 6242 8288
rect 7650 8236 7656 8288
rect 7708 8276 7714 8288
rect 7929 8279 7987 8285
rect 7929 8276 7941 8279
rect 7708 8248 7941 8276
rect 7708 8236 7714 8248
rect 7929 8245 7941 8248
rect 7975 8245 7987 8279
rect 7929 8239 7987 8245
rect 1104 8186 8280 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 8280 8186
rect 1104 8112 8280 8134
rect 3973 8075 4031 8081
rect 3973 8041 3985 8075
rect 4019 8072 4031 8075
rect 4062 8072 4068 8084
rect 4019 8044 4068 8072
rect 4019 8041 4031 8044
rect 3973 8035 4031 8041
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 5534 8032 5540 8084
rect 5592 8072 5598 8084
rect 6549 8075 6607 8081
rect 6549 8072 6561 8075
rect 5592 8044 6561 8072
rect 5592 8032 5598 8044
rect 6549 8041 6561 8044
rect 6595 8041 6607 8075
rect 6549 8035 6607 8041
rect 2961 8007 3019 8013
rect 2961 7973 2973 8007
rect 3007 8004 3019 8007
rect 3602 8004 3608 8016
rect 3007 7976 3608 8004
rect 3007 7973 3019 7976
rect 2961 7967 3019 7973
rect 3602 7964 3608 7976
rect 3660 7964 3666 8016
rect 3786 7964 3792 8016
rect 3844 8004 3850 8016
rect 4706 8004 4712 8016
rect 3844 7976 4712 8004
rect 3844 7964 3850 7976
rect 4706 7964 4712 7976
rect 4764 7964 4770 8016
rect 3510 7896 3516 7948
rect 3568 7936 3574 7948
rect 4062 7936 4068 7948
rect 3568 7908 4068 7936
rect 3568 7896 3574 7908
rect 4062 7896 4068 7908
rect 4120 7896 4126 7948
rect 4617 7939 4675 7945
rect 4617 7905 4629 7939
rect 4663 7936 4675 7939
rect 4890 7936 4896 7948
rect 4663 7908 4896 7936
rect 4663 7905 4675 7908
rect 4617 7899 4675 7905
rect 4890 7896 4896 7908
rect 4948 7936 4954 7948
rect 5258 7936 5264 7948
rect 4948 7908 5264 7936
rect 4948 7896 4954 7908
rect 5258 7896 5264 7908
rect 5316 7896 5322 7948
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7868 1639 7871
rect 2866 7868 2872 7880
rect 1627 7840 2872 7868
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 2866 7828 2872 7840
rect 2924 7828 2930 7880
rect 3145 7871 3203 7877
rect 3145 7837 3157 7871
rect 3191 7837 3203 7871
rect 3145 7831 3203 7837
rect 1848 7803 1906 7809
rect 1848 7769 1860 7803
rect 1894 7800 1906 7803
rect 2958 7800 2964 7812
rect 1894 7772 2964 7800
rect 1894 7769 1906 7772
rect 1848 7763 1906 7769
rect 2958 7760 2964 7772
rect 3016 7800 3022 7812
rect 3160 7800 3188 7831
rect 3602 7828 3608 7880
rect 3660 7828 3666 7880
rect 6362 7828 6368 7880
rect 6420 7868 6426 7880
rect 6457 7871 6515 7877
rect 6457 7868 6469 7871
rect 6420 7840 6469 7868
rect 6420 7828 6426 7840
rect 6457 7837 6469 7840
rect 6503 7868 6515 7871
rect 7929 7871 7987 7877
rect 7929 7868 7941 7871
rect 6503 7840 7941 7868
rect 6503 7837 6515 7840
rect 6457 7831 6515 7837
rect 7929 7837 7941 7840
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 3016 7772 3188 7800
rect 3016 7760 3022 7772
rect 4706 7760 4712 7812
rect 4764 7760 4770 7812
rect 7650 7800 7656 7812
rect 7708 7809 7714 7812
rect 7620 7772 7656 7800
rect 7650 7760 7656 7772
rect 7708 7763 7720 7809
rect 7708 7760 7714 7763
rect 1104 7642 8280 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 8280 7642
rect 1104 7568 8280 7590
rect 5353 7531 5411 7537
rect 5353 7497 5365 7531
rect 5399 7528 5411 7531
rect 5442 7528 5448 7540
rect 5399 7500 5448 7528
rect 5399 7497 5411 7500
rect 5353 7491 5411 7497
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 7466 7488 7472 7540
rect 7524 7528 7530 7540
rect 7745 7531 7803 7537
rect 7745 7528 7757 7531
rect 7524 7500 7757 7528
rect 7524 7488 7530 7500
rect 7745 7497 7757 7500
rect 7791 7497 7803 7531
rect 7745 7491 7803 7497
rect 2866 7460 2872 7472
rect 2516 7432 2872 7460
rect 2516 7401 2544 7432
rect 2866 7420 2872 7432
rect 2924 7460 2930 7472
rect 4240 7463 4298 7469
rect 2924 7432 4016 7460
rect 2924 7420 2930 7432
rect 2774 7401 2780 7404
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7361 2559 7395
rect 2501 7355 2559 7361
rect 2768 7355 2780 7401
rect 2774 7352 2780 7355
rect 2832 7352 2838 7404
rect 3988 7336 4016 7432
rect 4240 7429 4252 7463
rect 4286 7460 4298 7463
rect 4614 7460 4620 7472
rect 4286 7432 4620 7460
rect 4286 7429 4298 7432
rect 4240 7423 4298 7429
rect 4614 7420 4620 7432
rect 4672 7420 4678 7472
rect 6178 7420 6184 7472
rect 6236 7460 6242 7472
rect 6610 7463 6668 7469
rect 6610 7460 6622 7463
rect 6236 7432 6622 7460
rect 6236 7420 6242 7432
rect 6610 7429 6622 7432
rect 6656 7429 6668 7463
rect 6610 7423 6668 7429
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 5000 7364 5825 7392
rect 3970 7284 3976 7336
rect 4028 7284 4034 7336
rect 3418 7148 3424 7200
rect 3476 7188 3482 7200
rect 3881 7191 3939 7197
rect 3881 7188 3893 7191
rect 3476 7160 3893 7188
rect 3476 7148 3482 7160
rect 3881 7157 3893 7160
rect 3927 7188 3939 7191
rect 5000 7188 5028 7364
rect 5813 7361 5825 7364
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 6362 7352 6368 7404
rect 6420 7352 6426 7404
rect 5626 7284 5632 7336
rect 5684 7284 5690 7336
rect 5721 7327 5779 7333
rect 5721 7293 5733 7327
rect 5767 7324 5779 7327
rect 6270 7324 6276 7336
rect 5767 7296 6276 7324
rect 5767 7293 5779 7296
rect 5721 7287 5779 7293
rect 6270 7284 6276 7296
rect 6328 7284 6334 7336
rect 3927 7160 5028 7188
rect 3927 7157 3939 7160
rect 3881 7151 3939 7157
rect 6178 7148 6184 7200
rect 6236 7148 6242 7200
rect 1104 7098 8280 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 8280 7098
rect 1104 7024 8280 7046
rect 3896 6956 4936 6984
rect 3510 6916 3516 6928
rect 2148 6888 3516 6916
rect 2148 6860 2176 6888
rect 3510 6876 3516 6888
rect 3568 6876 3574 6928
rect 2130 6848 2136 6860
rect 2111 6820 2136 6848
rect 2130 6808 2136 6820
rect 2188 6808 2194 6860
rect 2682 6808 2688 6860
rect 2740 6848 2746 6860
rect 3896 6848 3924 6956
rect 2740 6820 3924 6848
rect 4908 6848 4936 6956
rect 5258 6944 5264 6996
rect 5316 6944 5322 6996
rect 5445 6851 5503 6857
rect 5445 6848 5457 6851
rect 4908 6820 5457 6848
rect 2740 6808 2746 6820
rect 5445 6817 5457 6820
rect 5491 6817 5503 6851
rect 5445 6811 5503 6817
rect 7098 6808 7104 6860
rect 7156 6848 7162 6860
rect 7745 6851 7803 6857
rect 7745 6848 7757 6851
rect 7156 6820 7757 6848
rect 7156 6808 7162 6820
rect 7745 6817 7757 6820
rect 7791 6817 7803 6851
rect 7745 6811 7803 6817
rect 1857 6783 1915 6789
rect 1857 6749 1869 6783
rect 1903 6749 1915 6783
rect 1857 6743 1915 6749
rect 1872 6712 1900 6743
rect 1946 6740 1952 6792
rect 2004 6740 2010 6792
rect 2314 6740 2320 6792
rect 2372 6740 2378 6792
rect 2590 6740 2596 6792
rect 2648 6780 2654 6792
rect 2961 6783 3019 6789
rect 2961 6780 2973 6783
rect 2648 6752 2973 6780
rect 2648 6740 2654 6752
rect 2961 6749 2973 6752
rect 3007 6749 3019 6783
rect 2961 6743 3019 6749
rect 3605 6783 3663 6789
rect 3605 6749 3617 6783
rect 3651 6780 3663 6783
rect 3786 6780 3792 6792
rect 3651 6752 3792 6780
rect 3651 6749 3663 6752
rect 3605 6743 3663 6749
rect 2869 6715 2927 6721
rect 1872 6684 2535 6712
rect 2133 6647 2191 6653
rect 2133 6613 2145 6647
rect 2179 6644 2191 6647
rect 2406 6644 2412 6656
rect 2179 6616 2412 6644
rect 2179 6613 2191 6616
rect 2133 6607 2191 6613
rect 2406 6604 2412 6616
rect 2464 6604 2470 6656
rect 2507 6644 2535 6684
rect 2869 6681 2881 6715
rect 2915 6712 2927 6715
rect 3050 6712 3056 6724
rect 2915 6684 3056 6712
rect 2915 6681 2927 6684
rect 2869 6675 2927 6681
rect 3050 6672 3056 6684
rect 3108 6672 3114 6724
rect 3620 6644 3648 6743
rect 3786 6740 3792 6752
rect 3844 6740 3850 6792
rect 3881 6783 3939 6789
rect 3881 6749 3893 6783
rect 3927 6780 3939 6783
rect 3970 6780 3976 6792
rect 3927 6752 3976 6780
rect 3927 6749 3939 6752
rect 3881 6743 3939 6749
rect 3970 6740 3976 6752
rect 4028 6780 4034 6792
rect 4028 6752 4292 6780
rect 4028 6740 4034 6752
rect 3694 6672 3700 6724
rect 3752 6712 3758 6724
rect 4126 6715 4184 6721
rect 4126 6712 4138 6715
rect 3752 6684 4138 6712
rect 3752 6672 3758 6684
rect 4126 6681 4138 6684
rect 4172 6681 4184 6715
rect 4264 6712 4292 6752
rect 4430 6740 4436 6792
rect 4488 6780 4494 6792
rect 5353 6783 5411 6789
rect 5353 6780 5365 6783
rect 4488 6752 5365 6780
rect 4488 6740 4494 6752
rect 5353 6749 5365 6752
rect 5399 6749 5411 6783
rect 5353 6743 5411 6749
rect 5534 6740 5540 6792
rect 5592 6740 5598 6792
rect 5721 6783 5779 6789
rect 5721 6749 5733 6783
rect 5767 6780 5779 6783
rect 6362 6780 6368 6792
rect 5767 6752 6368 6780
rect 5767 6749 5779 6752
rect 5721 6743 5779 6749
rect 5736 6712 5764 6743
rect 6362 6740 6368 6752
rect 6420 6740 6426 6792
rect 4264 6684 5764 6712
rect 5988 6715 6046 6721
rect 4126 6675 4184 6681
rect 5988 6681 6000 6715
rect 6034 6712 6046 6715
rect 6086 6712 6092 6724
rect 6034 6684 6092 6712
rect 6034 6681 6046 6684
rect 5988 6675 6046 6681
rect 6086 6672 6092 6684
rect 6144 6672 6150 6724
rect 2507 6616 3648 6644
rect 7098 6604 7104 6656
rect 7156 6604 7162 6656
rect 7193 6647 7251 6653
rect 7193 6613 7205 6647
rect 7239 6644 7251 6647
rect 7466 6644 7472 6656
rect 7239 6616 7472 6644
rect 7239 6613 7251 6616
rect 7193 6607 7251 6613
rect 7466 6604 7472 6616
rect 7524 6604 7530 6656
rect 7558 6604 7564 6656
rect 7616 6604 7622 6656
rect 7650 6604 7656 6656
rect 7708 6604 7714 6656
rect 1104 6554 8280 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 8280 6554
rect 1104 6480 8280 6502
rect 2590 6400 2596 6452
rect 2648 6400 2654 6452
rect 3878 6400 3884 6452
rect 3936 6440 3942 6452
rect 4249 6443 4307 6449
rect 4249 6440 4261 6443
rect 3936 6412 4261 6440
rect 3936 6400 3942 6412
rect 4249 6409 4261 6412
rect 4295 6409 4307 6443
rect 4249 6403 4307 6409
rect 4417 6443 4475 6449
rect 4417 6409 4429 6443
rect 4463 6440 4475 6443
rect 4890 6440 4896 6452
rect 4463 6412 4896 6440
rect 4463 6409 4475 6412
rect 4417 6403 4475 6409
rect 4890 6400 4896 6412
rect 4948 6440 4954 6452
rect 5350 6440 5356 6452
rect 4948 6412 5356 6440
rect 4948 6400 4954 6412
rect 5350 6400 5356 6412
rect 5408 6400 5414 6452
rect 6181 6443 6239 6449
rect 6181 6409 6193 6443
rect 6227 6440 6239 6443
rect 7650 6440 7656 6452
rect 6227 6412 7656 6440
rect 6227 6409 6239 6412
rect 6181 6403 6239 6409
rect 7650 6400 7656 6412
rect 7708 6400 7714 6452
rect 2406 6332 2412 6384
rect 2464 6332 2470 6384
rect 2866 6372 2872 6384
rect 2792 6344 2872 6372
rect 1946 6264 1952 6316
rect 2004 6304 2010 6316
rect 2685 6307 2743 6313
rect 2685 6304 2697 6307
rect 2004 6276 2697 6304
rect 2004 6264 2010 6276
rect 2685 6273 2697 6276
rect 2731 6304 2743 6307
rect 2792 6304 2820 6344
rect 2866 6332 2872 6344
rect 2924 6332 2930 6384
rect 3970 6372 3976 6384
rect 2976 6344 3976 6372
rect 2976 6304 3004 6344
rect 3970 6332 3976 6344
rect 4028 6332 4034 6384
rect 4617 6375 4675 6381
rect 4617 6341 4629 6375
rect 4663 6372 4675 6375
rect 7558 6372 7564 6384
rect 4663 6344 7564 6372
rect 4663 6341 4675 6344
rect 4617 6335 4675 6341
rect 3050 6313 3056 6316
rect 2731 6276 2820 6304
rect 2884 6276 3004 6304
rect 2731 6273 2743 6276
rect 2685 6267 2743 6273
rect 2777 6239 2835 6245
rect 2777 6205 2789 6239
rect 2823 6236 2835 6239
rect 2884 6236 2912 6276
rect 3044 6267 3056 6313
rect 3108 6304 3114 6316
rect 3108 6276 3144 6304
rect 3050 6264 3056 6267
rect 3108 6264 3114 6276
rect 2823 6208 2912 6236
rect 2823 6205 2835 6208
rect 2777 6199 2835 6205
rect 2314 6128 2320 6180
rect 2372 6168 2378 6180
rect 2409 6171 2467 6177
rect 2409 6168 2421 6171
rect 2372 6140 2421 6168
rect 2372 6128 2378 6140
rect 2409 6137 2421 6140
rect 2455 6137 2467 6171
rect 2409 6131 2467 6137
rect 3786 6128 3792 6180
rect 3844 6168 3850 6180
rect 4157 6171 4215 6177
rect 4157 6168 4169 6171
rect 3844 6140 4169 6168
rect 3844 6128 3850 6140
rect 4157 6137 4169 6140
rect 4203 6168 4215 6171
rect 4632 6168 4660 6335
rect 7558 6332 7564 6344
rect 7616 6332 7622 6384
rect 4982 6264 4988 6316
rect 5040 6304 5046 6316
rect 5169 6307 5227 6313
rect 5169 6304 5181 6307
rect 5040 6276 5181 6304
rect 5040 6264 5046 6276
rect 5169 6273 5181 6276
rect 5215 6273 5227 6307
rect 5169 6267 5227 6273
rect 6362 6264 6368 6316
rect 6420 6264 6426 6316
rect 6632 6307 6690 6313
rect 6632 6273 6644 6307
rect 6678 6304 6690 6307
rect 7190 6304 7196 6316
rect 6678 6276 7196 6304
rect 6678 6273 6690 6276
rect 6632 6267 6690 6273
rect 7190 6264 7196 6276
rect 7248 6264 7254 6316
rect 5077 6239 5135 6245
rect 5077 6205 5089 6239
rect 5123 6205 5135 6239
rect 5077 6199 5135 6205
rect 5261 6239 5319 6245
rect 5261 6205 5273 6239
rect 5307 6205 5319 6239
rect 5261 6199 5319 6205
rect 4203 6140 4660 6168
rect 4203 6137 4215 6140
rect 4157 6131 4215 6137
rect 3418 6060 3424 6112
rect 3476 6100 3482 6112
rect 4433 6103 4491 6109
rect 4433 6100 4445 6103
rect 3476 6072 4445 6100
rect 3476 6060 3482 6072
rect 4433 6069 4445 6072
rect 4479 6069 4491 6103
rect 4433 6063 4491 6069
rect 4798 6060 4804 6112
rect 4856 6100 4862 6112
rect 4893 6103 4951 6109
rect 4893 6100 4905 6103
rect 4856 6072 4905 6100
rect 4856 6060 4862 6072
rect 4893 6069 4905 6072
rect 4939 6069 4951 6103
rect 5092 6100 5120 6199
rect 5166 6128 5172 6180
rect 5224 6168 5230 6180
rect 5276 6168 5304 6199
rect 5350 6196 5356 6248
rect 5408 6196 5414 6248
rect 5629 6239 5687 6245
rect 5629 6205 5641 6239
rect 5675 6205 5687 6239
rect 5629 6199 5687 6205
rect 5224 6140 5304 6168
rect 5224 6128 5230 6140
rect 5258 6100 5264 6112
rect 5092 6072 5264 6100
rect 4893 6063 4951 6069
rect 5258 6060 5264 6072
rect 5316 6060 5322 6112
rect 5644 6100 5672 6199
rect 7650 6100 7656 6112
rect 5644 6072 7656 6100
rect 7650 6060 7656 6072
rect 7708 6100 7714 6112
rect 7745 6103 7803 6109
rect 7745 6100 7757 6103
rect 7708 6072 7757 6100
rect 7708 6060 7714 6072
rect 7745 6069 7757 6072
rect 7791 6069 7803 6103
rect 7745 6063 7803 6069
rect 1104 6010 8280 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 8280 6010
rect 1104 5936 8280 5958
rect 4706 5856 4712 5908
rect 4764 5896 4770 5908
rect 5353 5899 5411 5905
rect 5353 5896 5365 5899
rect 4764 5868 5365 5896
rect 4764 5856 4770 5868
rect 5353 5865 5365 5868
rect 5399 5865 5411 5899
rect 5353 5859 5411 5865
rect 6086 5856 6092 5908
rect 6144 5856 6150 5908
rect 6270 5856 6276 5908
rect 6328 5896 6334 5908
rect 6825 5899 6883 5905
rect 6825 5896 6837 5899
rect 6328 5868 6837 5896
rect 6328 5856 6334 5868
rect 6825 5865 6837 5868
rect 6871 5865 6883 5899
rect 6825 5859 6883 5865
rect 7834 5856 7840 5908
rect 7892 5856 7898 5908
rect 3605 5831 3663 5837
rect 3605 5797 3617 5831
rect 3651 5828 3663 5831
rect 5534 5828 5540 5840
rect 3651 5800 5540 5828
rect 3651 5797 3663 5800
rect 3605 5791 3663 5797
rect 5534 5788 5540 5800
rect 5592 5788 5598 5840
rect 2866 5720 2872 5772
rect 2924 5760 2930 5772
rect 4430 5760 4436 5772
rect 2924 5732 4436 5760
rect 2924 5720 2930 5732
rect 3160 5701 3188 5732
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 6178 5720 6184 5772
rect 6236 5760 6242 5772
rect 6641 5763 6699 5769
rect 6641 5760 6653 5763
rect 6236 5732 6653 5760
rect 6236 5720 6242 5732
rect 6641 5729 6653 5732
rect 6687 5729 6699 5763
rect 6641 5723 6699 5729
rect 7098 5720 7104 5772
rect 7156 5760 7162 5772
rect 7377 5763 7435 5769
rect 7377 5760 7389 5763
rect 7156 5732 7389 5760
rect 7156 5720 7162 5732
rect 7377 5729 7389 5732
rect 7423 5729 7435 5763
rect 7377 5723 7435 5729
rect 3145 5695 3203 5701
rect 3145 5661 3157 5695
rect 3191 5661 3203 5695
rect 3145 5655 3203 5661
rect 3418 5652 3424 5704
rect 3476 5652 3482 5704
rect 3694 5652 3700 5704
rect 3752 5692 3758 5704
rect 4982 5692 4988 5704
rect 3752 5664 4988 5692
rect 3752 5652 3758 5664
rect 4982 5652 4988 5664
rect 5040 5692 5046 5704
rect 5534 5692 5540 5704
rect 5040 5664 5540 5692
rect 5040 5652 5046 5664
rect 5534 5652 5540 5664
rect 5592 5652 5598 5704
rect 7392 5692 7420 5723
rect 7653 5695 7711 5701
rect 7653 5692 7665 5695
rect 7392 5664 7665 5692
rect 7653 5661 7665 5664
rect 7699 5661 7711 5695
rect 7653 5655 7711 5661
rect 3237 5627 3295 5633
rect 3237 5593 3249 5627
rect 3283 5624 3295 5627
rect 3786 5624 3792 5636
rect 3283 5596 3792 5624
rect 3283 5593 3295 5596
rect 3237 5587 3295 5593
rect 3786 5584 3792 5596
rect 3844 5584 3850 5636
rect 4062 5584 4068 5636
rect 4120 5584 4126 5636
rect 4430 5584 4436 5636
rect 4488 5624 4494 5636
rect 4890 5624 4896 5636
rect 4488 5596 4896 5624
rect 4488 5584 4494 5596
rect 4890 5584 4896 5596
rect 4948 5584 4954 5636
rect 3970 5516 3976 5568
rect 4028 5556 4034 5568
rect 5166 5556 5172 5568
rect 4028 5528 5172 5556
rect 4028 5516 4034 5528
rect 5166 5516 5172 5528
rect 5224 5516 5230 5568
rect 1104 5466 8280 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 8280 5466
rect 1104 5392 8280 5414
rect 4430 5312 4436 5364
rect 4488 5352 4494 5364
rect 4801 5355 4859 5361
rect 4801 5352 4813 5355
rect 4488 5324 4813 5352
rect 4488 5312 4494 5324
rect 4801 5321 4813 5324
rect 4847 5352 4859 5355
rect 4890 5352 4896 5364
rect 4847 5324 4896 5352
rect 4847 5321 4859 5324
rect 4801 5315 4859 5321
rect 4890 5312 4896 5324
rect 4948 5312 4954 5364
rect 4985 5355 5043 5361
rect 4985 5321 4997 5355
rect 5031 5352 5043 5355
rect 5350 5352 5356 5364
rect 5031 5324 5356 5352
rect 5031 5321 5043 5324
rect 4985 5315 5043 5321
rect 5350 5312 5356 5324
rect 5408 5352 5414 5364
rect 6733 5355 6791 5361
rect 6733 5352 6745 5355
rect 5408 5324 6745 5352
rect 5408 5312 5414 5324
rect 6733 5321 6745 5324
rect 6779 5321 6791 5355
rect 6733 5315 6791 5321
rect 7190 5312 7196 5364
rect 7248 5312 7254 5364
rect 2130 5244 2136 5296
rect 2188 5284 2194 5296
rect 2682 5284 2688 5296
rect 2188 5256 2688 5284
rect 2188 5244 2194 5256
rect 2682 5244 2688 5256
rect 2740 5244 2746 5296
rect 2901 5287 2959 5293
rect 2901 5253 2913 5287
rect 2947 5284 2959 5287
rect 4522 5284 4528 5296
rect 2947 5256 4528 5284
rect 2947 5253 2959 5256
rect 2901 5247 2959 5253
rect 4522 5244 4528 5256
rect 4580 5244 4586 5296
rect 5169 5287 5227 5293
rect 5169 5253 5181 5287
rect 5215 5253 5227 5287
rect 5169 5247 5227 5253
rect 3326 5176 3332 5228
rect 3384 5176 3390 5228
rect 4798 5216 4804 5228
rect 3436 5188 4804 5216
rect 3436 5148 3464 5188
rect 4798 5176 4804 5188
rect 4856 5176 4862 5228
rect 4982 5176 4988 5228
rect 5040 5216 5046 5228
rect 5077 5219 5135 5225
rect 5077 5216 5089 5219
rect 5040 5188 5089 5216
rect 5040 5176 5046 5188
rect 5077 5185 5089 5188
rect 5123 5185 5135 5219
rect 5184 5216 5212 5247
rect 5184 5188 5304 5216
rect 5077 5179 5135 5185
rect 2884 5120 3464 5148
rect 3605 5151 3663 5157
rect 2884 5021 2912 5120
rect 3605 5117 3617 5151
rect 3651 5148 3663 5151
rect 3970 5148 3976 5160
rect 3651 5120 3976 5148
rect 3651 5117 3663 5120
rect 3605 5111 3663 5117
rect 3970 5108 3976 5120
rect 4028 5108 4034 5160
rect 4065 5151 4123 5157
rect 4065 5117 4077 5151
rect 4111 5117 4123 5151
rect 5276 5148 5304 5188
rect 6086 5176 6092 5228
rect 6144 5216 6150 5228
rect 6825 5219 6883 5225
rect 6825 5216 6837 5219
rect 6144 5188 6837 5216
rect 6144 5176 6150 5188
rect 6825 5185 6837 5188
rect 6871 5185 6883 5219
rect 6825 5179 6883 5185
rect 7466 5176 7472 5228
rect 7524 5216 7530 5228
rect 7745 5219 7803 5225
rect 7745 5216 7757 5219
rect 7524 5188 7757 5216
rect 7524 5176 7530 5188
rect 7745 5185 7757 5188
rect 7791 5185 7803 5219
rect 7745 5179 7803 5185
rect 5534 5148 5540 5160
rect 5276 5120 5540 5148
rect 4065 5111 4123 5117
rect 3053 5083 3111 5089
rect 3053 5049 3065 5083
rect 3099 5080 3111 5083
rect 4080 5080 4108 5111
rect 5534 5108 5540 5120
rect 5592 5108 5598 5160
rect 5629 5151 5687 5157
rect 5629 5117 5641 5151
rect 5675 5117 5687 5151
rect 5629 5111 5687 5117
rect 5074 5080 5080 5092
rect 3099 5052 4016 5080
rect 4080 5052 5080 5080
rect 3099 5049 3111 5052
rect 3053 5043 3111 5049
rect 3988 5024 4016 5052
rect 5074 5040 5080 5052
rect 5132 5040 5138 5092
rect 5258 5040 5264 5092
rect 5316 5080 5322 5092
rect 5353 5083 5411 5089
rect 5353 5080 5365 5083
rect 5316 5052 5365 5080
rect 5316 5040 5322 5052
rect 5353 5049 5365 5052
rect 5399 5049 5411 5083
rect 5644 5080 5672 5111
rect 5994 5108 6000 5160
rect 6052 5148 6058 5160
rect 7006 5148 7012 5160
rect 6052 5120 7012 5148
rect 6052 5108 6058 5120
rect 7006 5108 7012 5120
rect 7064 5108 7070 5160
rect 6365 5083 6423 5089
rect 6365 5080 6377 5083
rect 5644 5052 6377 5080
rect 5353 5043 5411 5049
rect 6365 5049 6377 5052
rect 6411 5049 6423 5083
rect 6365 5043 6423 5049
rect 2869 5015 2927 5021
rect 2869 4981 2881 5015
rect 2915 4981 2927 5015
rect 2869 4975 2927 4981
rect 3142 4972 3148 5024
rect 3200 4972 3206 5024
rect 3513 5015 3571 5021
rect 3513 4981 3525 5015
rect 3559 5012 3571 5015
rect 3602 5012 3608 5024
rect 3559 4984 3608 5012
rect 3559 4981 3571 4984
rect 3513 4975 3571 4981
rect 3602 4972 3608 4984
rect 3660 4972 3666 5024
rect 3970 4972 3976 5024
rect 4028 4972 4034 5024
rect 4617 5015 4675 5021
rect 4617 4981 4629 5015
rect 4663 5012 4675 5015
rect 6086 5012 6092 5024
rect 4663 4984 6092 5012
rect 4663 4981 4675 4984
rect 4617 4975 4675 4981
rect 6086 4972 6092 4984
rect 6144 4972 6150 5024
rect 6178 4972 6184 5024
rect 6236 4972 6242 5024
rect 1104 4922 8280 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 8280 4922
rect 1104 4848 8280 4870
rect 3602 4768 3608 4820
rect 3660 4768 3666 4820
rect 3878 4768 3884 4820
rect 3936 4768 3942 4820
rect 5074 4768 5080 4820
rect 5132 4768 5138 4820
rect 5350 4768 5356 4820
rect 5408 4808 5414 4820
rect 5537 4811 5595 4817
rect 5537 4808 5549 4811
rect 5408 4780 5549 4808
rect 5408 4768 5414 4780
rect 5537 4777 5549 4780
rect 5583 4777 5595 4811
rect 7466 4808 7472 4820
rect 5537 4771 5595 4777
rect 6104 4780 7472 4808
rect 2593 4743 2651 4749
rect 2593 4709 2605 4743
rect 2639 4740 2651 4743
rect 2682 4740 2688 4752
rect 2639 4712 2688 4740
rect 2639 4709 2651 4712
rect 2593 4703 2651 4709
rect 2682 4700 2688 4712
rect 2740 4700 2746 4752
rect 3896 4740 3924 4768
rect 3804 4712 3924 4740
rect 5092 4740 5120 4768
rect 6104 4740 6132 4780
rect 7466 4768 7472 4780
rect 7524 4768 7530 4820
rect 7837 4811 7895 4817
rect 7837 4777 7849 4811
rect 7883 4808 7895 4811
rect 7926 4808 7932 4820
rect 7883 4780 7932 4808
rect 7883 4777 7895 4780
rect 7837 4771 7895 4777
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 5092 4712 6132 4740
rect 2869 4675 2927 4681
rect 2869 4641 2881 4675
rect 2915 4672 2927 4675
rect 3602 4672 3608 4684
rect 2915 4644 3608 4672
rect 2915 4641 2927 4644
rect 2869 4635 2927 4641
rect 3602 4632 3608 4644
rect 3660 4672 3666 4684
rect 3804 4672 3832 4712
rect 3660 4644 3832 4672
rect 3660 4632 3666 4644
rect 3804 4613 3832 4644
rect 3878 4632 3884 4684
rect 3936 4672 3942 4684
rect 4157 4675 4215 4681
rect 4157 4672 4169 4675
rect 3936 4644 4169 4672
rect 3936 4632 3942 4644
rect 4157 4641 4169 4644
rect 4203 4641 4215 4675
rect 4157 4635 4215 4641
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4573 3111 4607
rect 3053 4567 3111 4573
rect 3789 4607 3847 4613
rect 3789 4573 3801 4607
rect 3835 4573 3847 4607
rect 3789 4567 3847 4573
rect 3068 4536 3096 4567
rect 3970 4564 3976 4616
rect 4028 4604 4034 4616
rect 4413 4607 4471 4613
rect 4413 4604 4425 4607
rect 4028 4576 4425 4604
rect 4028 4564 4034 4576
rect 4413 4573 4425 4576
rect 4459 4573 4471 4607
rect 4413 4567 4471 4573
rect 5534 4564 5540 4616
rect 5592 4604 5598 4616
rect 5721 4607 5779 4613
rect 5721 4604 5733 4607
rect 5592 4576 5733 4604
rect 5592 4564 5598 4576
rect 5721 4573 5733 4576
rect 5767 4573 5779 4607
rect 5721 4567 5779 4573
rect 5810 4564 5816 4616
rect 5868 4604 5874 4616
rect 6089 4607 6147 4613
rect 6089 4604 6101 4607
rect 5868 4576 6101 4604
rect 5868 4564 5874 4576
rect 6089 4573 6101 4576
rect 6135 4573 6147 4607
rect 6089 4567 6147 4573
rect 6178 4564 6184 4616
rect 6236 4604 6242 4616
rect 6345 4607 6403 4613
rect 6345 4604 6357 4607
rect 6236 4576 6357 4604
rect 6236 4564 6242 4576
rect 6345 4573 6357 4576
rect 6391 4573 6403 4607
rect 6345 4567 6403 4573
rect 7650 4564 7656 4616
rect 7708 4564 7714 4616
rect 3234 4536 3240 4548
rect 3068 4508 3240 4536
rect 3234 4496 3240 4508
rect 3292 4536 3298 4548
rect 3694 4536 3700 4548
rect 3292 4508 3700 4536
rect 3292 4496 3298 4508
rect 3694 4496 3700 4508
rect 3752 4536 3758 4548
rect 3881 4539 3939 4545
rect 3881 4536 3893 4539
rect 3752 4508 3893 4536
rect 3752 4496 3758 4508
rect 3881 4505 3893 4508
rect 3927 4505 3939 4539
rect 3881 4499 3939 4505
rect 4065 4539 4123 4545
rect 4065 4505 4077 4539
rect 4111 4536 4123 4539
rect 4522 4536 4528 4548
rect 4111 4508 4528 4536
rect 4111 4505 4123 4508
rect 4065 4499 4123 4505
rect 4522 4496 4528 4508
rect 4580 4536 4586 4548
rect 4982 4536 4988 4548
rect 4580 4508 4988 4536
rect 4580 4496 4586 4508
rect 4982 4496 4988 4508
rect 5040 4496 5046 4548
rect 7742 4536 7748 4548
rect 5920 4508 7748 4536
rect 2406 4428 2412 4480
rect 2464 4428 2470 4480
rect 3786 4428 3792 4480
rect 3844 4428 3850 4480
rect 5920 4477 5948 4508
rect 7742 4496 7748 4508
rect 7800 4496 7806 4548
rect 5905 4471 5963 4477
rect 5905 4437 5917 4471
rect 5951 4437 5963 4471
rect 5905 4431 5963 4437
rect 1104 4378 8280 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 8280 4378
rect 1104 4304 8280 4326
rect 3694 4224 3700 4276
rect 3752 4264 3758 4276
rect 3789 4267 3847 4273
rect 3789 4264 3801 4267
rect 3752 4236 3801 4264
rect 3752 4224 3758 4236
rect 3789 4233 3801 4236
rect 3835 4233 3847 4267
rect 3789 4227 3847 4233
rect 4433 4199 4491 4205
rect 4433 4165 4445 4199
rect 4479 4196 4491 4199
rect 4706 4196 4712 4208
rect 4479 4168 4712 4196
rect 4479 4165 4491 4168
rect 4433 4159 4491 4165
rect 4706 4156 4712 4168
rect 4764 4156 4770 4208
rect 2676 4131 2734 4137
rect 2676 4097 2688 4131
rect 2722 4128 2734 4131
rect 3142 4128 3148 4140
rect 2722 4100 3148 4128
rect 2722 4097 2734 4100
rect 2676 4091 2734 4097
rect 3142 4088 3148 4100
rect 3200 4088 3206 4140
rect 4341 4131 4399 4137
rect 4341 4097 4353 4131
rect 4387 4128 4399 4131
rect 4798 4128 4804 4140
rect 4387 4100 4804 4128
rect 4387 4097 4399 4100
rect 4341 4091 4399 4097
rect 4798 4088 4804 4100
rect 4856 4088 4862 4140
rect 5350 4088 5356 4140
rect 5408 4128 5414 4140
rect 6621 4131 6679 4137
rect 6621 4128 6633 4131
rect 5408 4100 6633 4128
rect 5408 4088 5414 4100
rect 6621 4097 6633 4100
rect 6667 4097 6679 4131
rect 6621 4091 6679 4097
rect 2222 4020 2228 4072
rect 2280 4060 2286 4072
rect 2409 4063 2467 4069
rect 2409 4060 2421 4063
rect 2280 4032 2421 4060
rect 2280 4020 2286 4032
rect 2409 4029 2421 4032
rect 2455 4029 2467 4063
rect 2409 4023 2467 4029
rect 4249 4063 4307 4069
rect 4249 4029 4261 4063
rect 4295 4060 4307 4063
rect 4614 4060 4620 4072
rect 4295 4032 4620 4060
rect 4295 4029 4307 4032
rect 4249 4023 4307 4029
rect 4614 4020 4620 4032
rect 4672 4020 4678 4072
rect 5718 4020 5724 4072
rect 5776 4060 5782 4072
rect 6365 4063 6423 4069
rect 6365 4060 6377 4063
rect 5776 4032 6377 4060
rect 5776 4020 5782 4032
rect 6365 4029 6377 4032
rect 6411 4029 6423 4063
rect 6365 4023 6423 4029
rect 5718 3884 5724 3936
rect 5776 3884 5782 3936
rect 7650 3884 7656 3936
rect 7708 3924 7714 3936
rect 7745 3927 7803 3933
rect 7745 3924 7757 3927
rect 7708 3896 7757 3924
rect 7708 3884 7714 3896
rect 7745 3893 7757 3896
rect 7791 3893 7803 3927
rect 7745 3887 7803 3893
rect 1104 3834 8280 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 8280 3834
rect 1104 3760 8280 3782
rect 2222 3680 2228 3732
rect 2280 3720 2286 3732
rect 3878 3720 3884 3732
rect 2280 3692 3884 3720
rect 2280 3680 2286 3692
rect 3878 3680 3884 3692
rect 3936 3680 3942 3732
rect 4798 3680 4804 3732
rect 4856 3720 4862 3732
rect 5261 3723 5319 3729
rect 5261 3720 5273 3723
rect 4856 3692 5273 3720
rect 4856 3680 4862 3692
rect 5261 3689 5273 3692
rect 5307 3689 5319 3723
rect 5261 3683 5319 3689
rect 5534 3680 5540 3732
rect 5592 3720 5598 3732
rect 7377 3723 7435 3729
rect 7377 3720 7389 3723
rect 5592 3692 7389 3720
rect 5592 3680 5598 3692
rect 7377 3689 7389 3692
rect 7423 3689 7435 3723
rect 7377 3683 7435 3689
rect 7834 3680 7840 3732
rect 7892 3680 7898 3732
rect 3602 3612 3608 3664
rect 3660 3612 3666 3664
rect 2222 3544 2228 3596
rect 2280 3544 2286 3596
rect 3896 3593 3924 3680
rect 3881 3587 3939 3593
rect 3881 3553 3893 3587
rect 3927 3553 3939 3587
rect 3881 3547 3939 3553
rect 2492 3519 2550 3525
rect 2492 3485 2504 3519
rect 2538 3485 2550 3519
rect 3896 3516 3924 3547
rect 5445 3519 5503 3525
rect 5445 3516 5457 3519
rect 3896 3488 5457 3516
rect 2492 3479 2550 3485
rect 5445 3485 5457 3488
rect 5491 3516 5503 3519
rect 5718 3516 5724 3528
rect 5491 3488 5724 3516
rect 5491 3485 5503 3488
rect 5445 3479 5503 3485
rect 2406 3408 2412 3460
rect 2464 3448 2470 3460
rect 2516 3448 2544 3479
rect 5718 3476 5724 3488
rect 5776 3516 5782 3528
rect 5997 3519 6055 3525
rect 5997 3516 6009 3519
rect 5776 3488 6009 3516
rect 5776 3476 5782 3488
rect 5997 3485 6009 3488
rect 6043 3516 6055 3519
rect 6086 3516 6092 3528
rect 6043 3488 6092 3516
rect 6043 3485 6055 3488
rect 5997 3479 6055 3485
rect 6086 3476 6092 3488
rect 6144 3476 6150 3528
rect 7466 3476 7472 3528
rect 7524 3516 7530 3528
rect 7653 3519 7711 3525
rect 7653 3516 7665 3519
rect 7524 3488 7665 3516
rect 7524 3476 7530 3488
rect 7653 3485 7665 3488
rect 7699 3485 7711 3519
rect 7653 3479 7711 3485
rect 2464 3420 2544 3448
rect 2464 3408 2470 3420
rect 3694 3408 3700 3460
rect 3752 3448 3758 3460
rect 4126 3451 4184 3457
rect 4126 3448 4138 3451
rect 3752 3420 4138 3448
rect 3752 3408 3758 3420
rect 4126 3417 4138 3420
rect 4172 3417 4184 3451
rect 4126 3411 4184 3417
rect 5902 3408 5908 3460
rect 5960 3448 5966 3460
rect 6242 3451 6300 3457
rect 6242 3448 6254 3451
rect 5960 3420 6254 3448
rect 5960 3408 5966 3420
rect 6242 3417 6254 3420
rect 6288 3417 6300 3451
rect 6242 3411 6300 3417
rect 4338 3340 4344 3392
rect 4396 3380 4402 3392
rect 7650 3380 7656 3392
rect 4396 3352 7656 3380
rect 4396 3340 4402 3352
rect 7650 3340 7656 3352
rect 7708 3340 7714 3392
rect 1104 3290 8280 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 8280 3290
rect 1104 3216 8280 3238
rect 2961 3179 3019 3185
rect 2961 3145 2973 3179
rect 3007 3176 3019 3179
rect 3326 3176 3332 3188
rect 3007 3148 3332 3176
rect 3007 3145 3019 3148
rect 2961 3139 3019 3145
rect 3326 3136 3332 3148
rect 3384 3136 3390 3188
rect 5350 3136 5356 3188
rect 5408 3136 5414 3188
rect 7745 3179 7803 3185
rect 7745 3145 7757 3179
rect 7791 3145 7803 3179
rect 7745 3139 7803 3145
rect 4617 3111 4675 3117
rect 4617 3077 4629 3111
rect 4663 3108 4675 3111
rect 5905 3111 5963 3117
rect 5905 3108 5917 3111
rect 4663 3080 5917 3108
rect 4663 3077 4675 3080
rect 4617 3071 4675 3077
rect 5905 3077 5917 3080
rect 5951 3077 5963 3111
rect 7760 3108 7788 3139
rect 5905 3071 5963 3077
rect 6012 3080 7788 3108
rect 3053 3043 3111 3049
rect 3053 3009 3065 3043
rect 3099 3009 3111 3043
rect 3053 3003 3111 3009
rect 3145 3043 3203 3049
rect 3145 3009 3157 3043
rect 3191 3040 3203 3043
rect 3234 3040 3240 3052
rect 3191 3012 3240 3040
rect 3191 3009 3203 3012
rect 3145 3003 3203 3009
rect 2682 2932 2688 2984
rect 2740 2932 2746 2984
rect 3068 2972 3096 3003
rect 3234 3000 3240 3012
rect 3292 3000 3298 3052
rect 3326 3000 3332 3052
rect 3384 3040 3390 3052
rect 3384 3012 4936 3040
rect 3384 3000 3390 3012
rect 3602 2972 3608 2984
rect 3068 2944 3608 2972
rect 3602 2932 3608 2944
rect 3660 2972 3666 2984
rect 3970 2972 3976 2984
rect 3660 2944 3976 2972
rect 3660 2932 3666 2944
rect 3970 2932 3976 2944
rect 4028 2932 4034 2984
rect 4065 2975 4123 2981
rect 4065 2941 4077 2975
rect 4111 2972 4123 2975
rect 4338 2972 4344 2984
rect 4111 2944 4344 2972
rect 4111 2941 4123 2944
rect 4065 2935 4123 2941
rect 4338 2932 4344 2944
rect 4396 2932 4402 2984
rect 4801 2975 4859 2981
rect 4801 2941 4813 2975
rect 4847 2941 4859 2975
rect 4908 2972 4936 3012
rect 4982 3000 4988 3052
rect 5040 3040 5046 3052
rect 5813 3043 5871 3049
rect 5813 3040 5825 3043
rect 5040 3012 5825 3040
rect 5040 3000 5046 3012
rect 5813 3009 5825 3012
rect 5859 3009 5871 3043
rect 6012 3040 6040 3080
rect 5813 3003 5871 3009
rect 5920 3012 6040 3040
rect 5920 2972 5948 3012
rect 6086 3000 6092 3052
rect 6144 3040 6150 3052
rect 6638 3049 6644 3052
rect 6365 3043 6423 3049
rect 6365 3040 6377 3043
rect 6144 3012 6377 3040
rect 6144 3000 6150 3012
rect 6365 3009 6377 3012
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 6632 3003 6644 3049
rect 6638 3000 6644 3003
rect 6696 3000 6702 3052
rect 4908 2944 5948 2972
rect 4801 2935 4859 2941
rect 4816 2904 4844 2935
rect 5994 2932 6000 2984
rect 6052 2932 6058 2984
rect 5445 2907 5503 2913
rect 5445 2904 5457 2907
rect 4816 2876 5457 2904
rect 5445 2873 5457 2876
rect 5491 2873 5503 2907
rect 5445 2867 5503 2873
rect 3881 2839 3939 2845
rect 3881 2805 3893 2839
rect 3927 2836 3939 2839
rect 7098 2836 7104 2848
rect 3927 2808 7104 2836
rect 3927 2805 3939 2808
rect 3881 2799 3939 2805
rect 7098 2796 7104 2808
rect 7156 2796 7162 2848
rect 1104 2746 8280 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 8280 2746
rect 1104 2672 8280 2694
rect 3421 2635 3479 2641
rect 3421 2601 3433 2635
rect 3467 2632 3479 2635
rect 3881 2635 3939 2641
rect 3881 2632 3893 2635
rect 3467 2604 3893 2632
rect 3467 2601 3479 2604
rect 3421 2595 3479 2601
rect 3881 2601 3893 2604
rect 3927 2601 3939 2635
rect 3881 2595 3939 2601
rect 5902 2592 5908 2644
rect 5960 2592 5966 2644
rect 6638 2592 6644 2644
rect 6696 2592 6702 2644
rect 7834 2592 7840 2644
rect 7892 2592 7898 2644
rect 3605 2567 3663 2573
rect 3605 2533 3617 2567
rect 3651 2564 3663 2567
rect 3694 2564 3700 2576
rect 3651 2536 3700 2564
rect 3651 2533 3663 2536
rect 3605 2527 3663 2533
rect 3694 2524 3700 2536
rect 3752 2524 3758 2576
rect 4890 2524 4896 2576
rect 4948 2564 4954 2576
rect 5258 2564 5264 2576
rect 4948 2536 5264 2564
rect 4948 2524 4954 2536
rect 5258 2524 5264 2536
rect 5316 2564 5322 2576
rect 5316 2536 7328 2564
rect 5316 2524 5322 2536
rect 3234 2456 3240 2508
rect 3292 2496 3298 2508
rect 4798 2496 4804 2508
rect 3292 2468 4016 2496
rect 3292 2456 3298 2468
rect 3145 2431 3203 2437
rect 3145 2397 3157 2431
rect 3191 2428 3203 2431
rect 3326 2428 3332 2440
rect 3191 2400 3332 2428
rect 3191 2397 3203 2400
rect 3145 2391 3203 2397
rect 3326 2388 3332 2400
rect 3384 2388 3390 2440
rect 2682 2320 2688 2372
rect 2740 2360 2746 2372
rect 3237 2363 3295 2369
rect 3237 2360 3249 2363
rect 2740 2332 3249 2360
rect 2740 2320 2746 2332
rect 3237 2329 3249 2332
rect 3283 2329 3295 2363
rect 3237 2323 3295 2329
rect 3453 2363 3511 2369
rect 3453 2329 3465 2363
rect 3499 2360 3511 2363
rect 3786 2360 3792 2372
rect 3499 2332 3792 2360
rect 3499 2329 3511 2332
rect 3453 2323 3511 2329
rect 3786 2320 3792 2332
rect 3844 2320 3850 2372
rect 3988 2360 4016 2468
rect 4080 2468 4804 2496
rect 4080 2437 4108 2468
rect 4798 2456 4804 2468
rect 4856 2456 4862 2508
rect 5353 2499 5411 2505
rect 5353 2465 5365 2499
rect 5399 2496 5411 2499
rect 5994 2496 6000 2508
rect 5399 2468 6000 2496
rect 5399 2465 5411 2468
rect 5353 2459 5411 2465
rect 5994 2456 6000 2468
rect 6052 2456 6058 2508
rect 7098 2456 7104 2508
rect 7156 2456 7162 2508
rect 7193 2499 7251 2505
rect 7193 2465 7205 2499
rect 7239 2465 7251 2499
rect 7193 2459 7251 2465
rect 4065 2431 4123 2437
rect 4065 2397 4077 2431
rect 4111 2397 4123 2431
rect 4065 2391 4123 2397
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2397 4399 2431
rect 4341 2391 4399 2397
rect 4525 2431 4583 2437
rect 4525 2397 4537 2431
rect 4571 2428 4583 2431
rect 5534 2428 5540 2440
rect 4571 2400 5540 2428
rect 4571 2397 4583 2400
rect 4525 2391 4583 2397
rect 4356 2360 4384 2391
rect 5534 2388 5540 2400
rect 5592 2388 5598 2440
rect 6012 2428 6040 2456
rect 7208 2428 7236 2459
rect 6012 2400 7236 2428
rect 7009 2363 7067 2369
rect 3988 2332 5580 2360
rect 2958 2252 2964 2304
rect 3016 2252 3022 2304
rect 4154 2252 4160 2304
rect 4212 2292 4218 2304
rect 4249 2295 4307 2301
rect 4249 2292 4261 2295
rect 4212 2264 4261 2292
rect 4212 2252 4218 2264
rect 4249 2261 4261 2264
rect 4295 2292 4307 2295
rect 4890 2292 4896 2304
rect 4295 2264 4896 2292
rect 4295 2261 4307 2264
rect 4249 2255 4307 2261
rect 4890 2252 4896 2264
rect 4948 2252 4954 2304
rect 5552 2301 5580 2332
rect 7009 2329 7021 2363
rect 7055 2360 7067 2363
rect 7300 2360 7328 2536
rect 7650 2388 7656 2440
rect 7708 2388 7714 2440
rect 7055 2332 7328 2360
rect 7055 2329 7067 2332
rect 7009 2323 7067 2329
rect 5077 2295 5135 2301
rect 5077 2261 5089 2295
rect 5123 2292 5135 2295
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 5123 2264 5457 2292
rect 5123 2261 5135 2264
rect 5077 2255 5135 2261
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 5445 2255 5503 2261
rect 5537 2295 5595 2301
rect 5537 2261 5549 2295
rect 5583 2261 5595 2295
rect 5537 2255 5595 2261
rect 1104 2202 8280 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 8280 2202
rect 1104 2128 8280 2150
rect 2958 2048 2964 2100
rect 3016 2088 3022 2100
rect 6914 2088 6920 2100
rect 3016 2060 6920 2088
rect 3016 2048 3022 2060
rect 6914 2048 6920 2060
rect 6972 2048 6978 2100
<< via1 >>
rect 3056 9324 3108 9376
rect 5540 9324 5592 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 6920 9120 6972 9172
rect 7656 9163 7708 9172
rect 7656 9129 7665 9163
rect 7665 9129 7699 9163
rect 7699 9129 7708 9163
rect 7656 9120 7708 9129
rect 848 8916 900 8968
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 3424 8916 3476 8968
rect 3700 8984 3752 9036
rect 3792 8916 3844 8968
rect 4068 8959 4120 8968
rect 4068 8925 4077 8959
rect 4077 8925 4111 8959
rect 4111 8925 4120 8959
rect 4068 8916 4120 8925
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4160 8916 4212 8925
rect 5448 8984 5500 9036
rect 2964 8848 3016 8900
rect 5264 8916 5316 8968
rect 5540 8959 5592 8968
rect 5540 8925 5549 8959
rect 5549 8925 5583 8959
rect 5583 8925 5592 8959
rect 5540 8916 5592 8925
rect 7104 8984 7156 9036
rect 7472 8959 7524 8968
rect 7472 8925 7481 8959
rect 7481 8925 7515 8959
rect 7515 8925 7524 8959
rect 7472 8916 7524 8925
rect 3976 8780 4028 8832
rect 4620 8780 4672 8832
rect 6184 8823 6236 8832
rect 6184 8789 6193 8823
rect 6193 8789 6227 8823
rect 6227 8789 6236 8823
rect 6184 8780 6236 8789
rect 6644 8823 6696 8832
rect 6644 8789 6653 8823
rect 6653 8789 6687 8823
rect 6687 8789 6696 8823
rect 6644 8780 6696 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 3700 8576 3752 8628
rect 3792 8576 3844 8628
rect 2688 8483 2740 8492
rect 2688 8449 2697 8483
rect 2697 8449 2731 8483
rect 2731 8449 2740 8483
rect 2688 8440 2740 8449
rect 2964 8483 3016 8492
rect 2964 8449 2973 8483
rect 2973 8449 3007 8483
rect 3007 8449 3016 8483
rect 2964 8440 3016 8449
rect 3608 8440 3660 8492
rect 4896 8508 4948 8560
rect 6184 8576 6236 8628
rect 3976 8483 4028 8492
rect 3976 8449 3985 8483
rect 3985 8449 4019 8483
rect 4019 8449 4028 8483
rect 3976 8440 4028 8449
rect 4252 8483 4304 8492
rect 4252 8449 4261 8483
rect 4261 8449 4295 8483
rect 4295 8449 4304 8483
rect 4252 8440 4304 8449
rect 4436 8483 4488 8492
rect 4436 8449 4445 8483
rect 4445 8449 4479 8483
rect 4479 8449 4488 8483
rect 4436 8440 4488 8449
rect 4712 8440 4764 8492
rect 5264 8440 5316 8492
rect 5448 8483 5500 8492
rect 5448 8449 5457 8483
rect 5457 8449 5491 8483
rect 5491 8449 5500 8483
rect 5448 8440 5500 8449
rect 6644 8440 6696 8492
rect 2780 8304 2832 8356
rect 3700 8304 3752 8356
rect 4252 8304 4304 8356
rect 5356 8304 5408 8356
rect 7104 8372 7156 8424
rect 5632 8236 5684 8288
rect 6184 8279 6236 8288
rect 6184 8245 6193 8279
rect 6193 8245 6227 8279
rect 6227 8245 6236 8279
rect 6184 8236 6236 8245
rect 7656 8236 7708 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 4068 8032 4120 8084
rect 5540 8032 5592 8084
rect 3608 7964 3660 8016
rect 3792 7964 3844 8016
rect 4712 7964 4764 8016
rect 3516 7939 3568 7948
rect 3516 7905 3525 7939
rect 3525 7905 3559 7939
rect 3559 7905 3568 7939
rect 3516 7896 3568 7905
rect 4068 7896 4120 7948
rect 4896 7896 4948 7948
rect 5264 7896 5316 7948
rect 2872 7828 2924 7880
rect 2964 7760 3016 7812
rect 3608 7871 3660 7880
rect 3608 7837 3617 7871
rect 3617 7837 3651 7871
rect 3651 7837 3660 7871
rect 3608 7828 3660 7837
rect 6368 7828 6420 7880
rect 4712 7803 4764 7812
rect 4712 7769 4721 7803
rect 4721 7769 4755 7803
rect 4755 7769 4764 7803
rect 4712 7760 4764 7769
rect 7656 7803 7708 7812
rect 7656 7769 7674 7803
rect 7674 7769 7708 7803
rect 7656 7760 7708 7769
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 5448 7488 5500 7540
rect 7472 7488 7524 7540
rect 2872 7420 2924 7472
rect 2780 7395 2832 7404
rect 2780 7361 2814 7395
rect 2814 7361 2832 7395
rect 2780 7352 2832 7361
rect 4620 7420 4672 7472
rect 6184 7420 6236 7472
rect 3976 7327 4028 7336
rect 3976 7293 3985 7327
rect 3985 7293 4019 7327
rect 4019 7293 4028 7327
rect 3976 7284 4028 7293
rect 3424 7148 3476 7200
rect 6368 7395 6420 7404
rect 6368 7361 6377 7395
rect 6377 7361 6411 7395
rect 6411 7361 6420 7395
rect 6368 7352 6420 7361
rect 5632 7327 5684 7336
rect 5632 7293 5641 7327
rect 5641 7293 5675 7327
rect 5675 7293 5684 7327
rect 5632 7284 5684 7293
rect 6276 7284 6328 7336
rect 6184 7191 6236 7200
rect 6184 7157 6193 7191
rect 6193 7157 6227 7191
rect 6227 7157 6236 7191
rect 6184 7148 6236 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 3516 6876 3568 6928
rect 2136 6851 2188 6860
rect 2136 6817 2145 6851
rect 2145 6817 2179 6851
rect 2179 6817 2188 6851
rect 2136 6808 2188 6817
rect 2688 6808 2740 6860
rect 5264 6987 5316 6996
rect 5264 6953 5273 6987
rect 5273 6953 5307 6987
rect 5307 6953 5316 6987
rect 5264 6944 5316 6953
rect 7104 6808 7156 6860
rect 1952 6783 2004 6792
rect 1952 6749 1961 6783
rect 1961 6749 1995 6783
rect 1995 6749 2004 6783
rect 1952 6740 2004 6749
rect 2320 6783 2372 6792
rect 2320 6749 2329 6783
rect 2329 6749 2363 6783
rect 2363 6749 2372 6783
rect 2320 6740 2372 6749
rect 2596 6740 2648 6792
rect 2412 6604 2464 6656
rect 3056 6672 3108 6724
rect 3792 6740 3844 6792
rect 3976 6740 4028 6792
rect 3700 6672 3752 6724
rect 4436 6740 4488 6792
rect 5540 6783 5592 6792
rect 5540 6749 5549 6783
rect 5549 6749 5583 6783
rect 5583 6749 5592 6783
rect 5540 6740 5592 6749
rect 6368 6740 6420 6792
rect 6092 6672 6144 6724
rect 7104 6647 7156 6656
rect 7104 6613 7113 6647
rect 7113 6613 7147 6647
rect 7147 6613 7156 6647
rect 7104 6604 7156 6613
rect 7472 6604 7524 6656
rect 7564 6647 7616 6656
rect 7564 6613 7573 6647
rect 7573 6613 7607 6647
rect 7607 6613 7616 6647
rect 7564 6604 7616 6613
rect 7656 6647 7708 6656
rect 7656 6613 7665 6647
rect 7665 6613 7699 6647
rect 7699 6613 7708 6647
rect 7656 6604 7708 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 2596 6443 2648 6452
rect 2596 6409 2605 6443
rect 2605 6409 2639 6443
rect 2639 6409 2648 6443
rect 2596 6400 2648 6409
rect 3884 6400 3936 6452
rect 4896 6400 4948 6452
rect 5356 6400 5408 6452
rect 7656 6400 7708 6452
rect 2412 6375 2464 6384
rect 2412 6341 2421 6375
rect 2421 6341 2455 6375
rect 2455 6341 2464 6375
rect 2412 6332 2464 6341
rect 1952 6264 2004 6316
rect 2872 6332 2924 6384
rect 3976 6332 4028 6384
rect 3056 6307 3108 6316
rect 3056 6273 3090 6307
rect 3090 6273 3108 6307
rect 3056 6264 3108 6273
rect 2320 6128 2372 6180
rect 3792 6128 3844 6180
rect 7564 6332 7616 6384
rect 4988 6264 5040 6316
rect 6368 6307 6420 6316
rect 6368 6273 6377 6307
rect 6377 6273 6411 6307
rect 6411 6273 6420 6307
rect 6368 6264 6420 6273
rect 7196 6264 7248 6316
rect 3424 6060 3476 6112
rect 4804 6060 4856 6112
rect 5172 6128 5224 6180
rect 5356 6239 5408 6248
rect 5356 6205 5365 6239
rect 5365 6205 5399 6239
rect 5399 6205 5408 6239
rect 5356 6196 5408 6205
rect 5264 6060 5316 6112
rect 7656 6060 7708 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 4712 5856 4764 5908
rect 6092 5899 6144 5908
rect 6092 5865 6101 5899
rect 6101 5865 6135 5899
rect 6135 5865 6144 5899
rect 6092 5856 6144 5865
rect 6276 5856 6328 5908
rect 7840 5899 7892 5908
rect 7840 5865 7849 5899
rect 7849 5865 7883 5899
rect 7883 5865 7892 5899
rect 7840 5856 7892 5865
rect 5540 5788 5592 5840
rect 2872 5720 2924 5772
rect 4436 5720 4488 5772
rect 6184 5720 6236 5772
rect 7104 5720 7156 5772
rect 3424 5695 3476 5704
rect 3424 5661 3433 5695
rect 3433 5661 3467 5695
rect 3467 5661 3476 5695
rect 3424 5652 3476 5661
rect 3700 5652 3752 5704
rect 4988 5652 5040 5704
rect 5540 5652 5592 5704
rect 3792 5584 3844 5636
rect 4068 5627 4120 5636
rect 4068 5593 4077 5627
rect 4077 5593 4111 5627
rect 4111 5593 4120 5627
rect 4068 5584 4120 5593
rect 4436 5584 4488 5636
rect 4896 5584 4948 5636
rect 3976 5516 4028 5568
rect 5172 5516 5224 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 4436 5312 4488 5364
rect 4896 5312 4948 5364
rect 5356 5312 5408 5364
rect 7196 5355 7248 5364
rect 7196 5321 7205 5355
rect 7205 5321 7239 5355
rect 7239 5321 7248 5355
rect 7196 5312 7248 5321
rect 2136 5244 2188 5296
rect 2688 5287 2740 5296
rect 2688 5253 2697 5287
rect 2697 5253 2731 5287
rect 2731 5253 2740 5287
rect 2688 5244 2740 5253
rect 4528 5244 4580 5296
rect 3332 5219 3384 5228
rect 3332 5185 3341 5219
rect 3341 5185 3375 5219
rect 3375 5185 3384 5219
rect 3332 5176 3384 5185
rect 4804 5176 4856 5228
rect 4988 5176 5040 5228
rect 3976 5108 4028 5160
rect 6092 5176 6144 5228
rect 7472 5176 7524 5228
rect 5540 5108 5592 5160
rect 5080 5040 5132 5092
rect 5264 5040 5316 5092
rect 6000 5108 6052 5160
rect 7012 5151 7064 5160
rect 7012 5117 7021 5151
rect 7021 5117 7055 5151
rect 7055 5117 7064 5151
rect 7012 5108 7064 5117
rect 3148 5015 3200 5024
rect 3148 4981 3157 5015
rect 3157 4981 3191 5015
rect 3191 4981 3200 5015
rect 3148 4972 3200 4981
rect 3608 4972 3660 5024
rect 3976 4972 4028 5024
rect 6092 4972 6144 5024
rect 6184 5015 6236 5024
rect 6184 4981 6193 5015
rect 6193 4981 6227 5015
rect 6227 4981 6236 5015
rect 6184 4972 6236 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 3608 4811 3660 4820
rect 3608 4777 3617 4811
rect 3617 4777 3651 4811
rect 3651 4777 3660 4811
rect 3608 4768 3660 4777
rect 3884 4768 3936 4820
rect 5080 4768 5132 4820
rect 5356 4768 5408 4820
rect 7472 4811 7524 4820
rect 2688 4700 2740 4752
rect 7472 4777 7481 4811
rect 7481 4777 7515 4811
rect 7515 4777 7524 4811
rect 7472 4768 7524 4777
rect 7932 4768 7984 4820
rect 3608 4632 3660 4684
rect 3884 4632 3936 4684
rect 3976 4564 4028 4616
rect 5540 4564 5592 4616
rect 5816 4564 5868 4616
rect 6184 4564 6236 4616
rect 7656 4607 7708 4616
rect 7656 4573 7665 4607
rect 7665 4573 7699 4607
rect 7699 4573 7708 4607
rect 7656 4564 7708 4573
rect 3240 4496 3292 4548
rect 3700 4496 3752 4548
rect 4528 4496 4580 4548
rect 4988 4496 5040 4548
rect 2412 4471 2464 4480
rect 2412 4437 2421 4471
rect 2421 4437 2455 4471
rect 2455 4437 2464 4471
rect 2412 4428 2464 4437
rect 3792 4471 3844 4480
rect 3792 4437 3801 4471
rect 3801 4437 3835 4471
rect 3835 4437 3844 4471
rect 3792 4428 3844 4437
rect 7748 4496 7800 4548
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 3700 4224 3752 4276
rect 4712 4156 4764 4208
rect 3148 4088 3200 4140
rect 4804 4088 4856 4140
rect 5356 4088 5408 4140
rect 2228 4020 2280 4072
rect 4620 4020 4672 4072
rect 5724 4020 5776 4072
rect 5724 3927 5776 3936
rect 5724 3893 5733 3927
rect 5733 3893 5767 3927
rect 5767 3893 5776 3927
rect 5724 3884 5776 3893
rect 7656 3884 7708 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 2228 3680 2280 3732
rect 3884 3680 3936 3732
rect 4804 3680 4856 3732
rect 5540 3680 5592 3732
rect 7840 3723 7892 3732
rect 7840 3689 7849 3723
rect 7849 3689 7883 3723
rect 7883 3689 7892 3723
rect 7840 3680 7892 3689
rect 3608 3655 3660 3664
rect 3608 3621 3617 3655
rect 3617 3621 3651 3655
rect 3651 3621 3660 3655
rect 3608 3612 3660 3621
rect 2228 3587 2280 3596
rect 2228 3553 2237 3587
rect 2237 3553 2271 3587
rect 2271 3553 2280 3587
rect 2228 3544 2280 3553
rect 2412 3408 2464 3460
rect 5724 3476 5776 3528
rect 6092 3476 6144 3528
rect 7472 3476 7524 3528
rect 3700 3408 3752 3460
rect 5908 3408 5960 3460
rect 4344 3340 4396 3392
rect 7656 3340 7708 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 3332 3136 3384 3188
rect 5356 3179 5408 3188
rect 5356 3145 5365 3179
rect 5365 3145 5399 3179
rect 5399 3145 5408 3179
rect 5356 3136 5408 3145
rect 2688 2975 2740 2984
rect 2688 2941 2697 2975
rect 2697 2941 2731 2975
rect 2731 2941 2740 2975
rect 2688 2932 2740 2941
rect 3240 3000 3292 3052
rect 3332 3043 3384 3052
rect 3332 3009 3341 3043
rect 3341 3009 3375 3043
rect 3375 3009 3384 3043
rect 3332 3000 3384 3009
rect 3608 2932 3660 2984
rect 3976 2932 4028 2984
rect 4344 2932 4396 2984
rect 4988 3000 5040 3052
rect 6092 3000 6144 3052
rect 6644 3043 6696 3052
rect 6644 3009 6678 3043
rect 6678 3009 6696 3043
rect 6644 3000 6696 3009
rect 6000 2975 6052 2984
rect 6000 2941 6009 2975
rect 6009 2941 6043 2975
rect 6043 2941 6052 2975
rect 6000 2932 6052 2941
rect 7104 2796 7156 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 5908 2635 5960 2644
rect 5908 2601 5917 2635
rect 5917 2601 5951 2635
rect 5951 2601 5960 2635
rect 5908 2592 5960 2601
rect 6644 2635 6696 2644
rect 6644 2601 6653 2635
rect 6653 2601 6687 2635
rect 6687 2601 6696 2635
rect 6644 2592 6696 2601
rect 7840 2635 7892 2644
rect 7840 2601 7849 2635
rect 7849 2601 7883 2635
rect 7883 2601 7892 2635
rect 7840 2592 7892 2601
rect 3700 2524 3752 2576
rect 4896 2524 4948 2576
rect 5264 2524 5316 2576
rect 3240 2456 3292 2508
rect 3332 2388 3384 2440
rect 2688 2320 2740 2372
rect 3792 2320 3844 2372
rect 4804 2456 4856 2508
rect 6000 2456 6052 2508
rect 7104 2499 7156 2508
rect 7104 2465 7113 2499
rect 7113 2465 7147 2499
rect 7147 2465 7156 2499
rect 7104 2456 7156 2465
rect 5540 2388 5592 2440
rect 2964 2295 3016 2304
rect 2964 2261 2973 2295
rect 2973 2261 3007 2295
rect 3007 2261 3016 2295
rect 2964 2252 3016 2261
rect 4160 2252 4212 2304
rect 4896 2252 4948 2304
rect 7656 2431 7708 2440
rect 7656 2397 7665 2431
rect 7665 2397 7699 2431
rect 7699 2397 7708 2431
rect 7656 2388 7708 2397
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 2964 2048 3016 2100
rect 6920 2048 6972 2100
<< metal2 >>
rect 7654 10432 7710 10441
rect 7654 10367 7710 10376
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 3068 8974 3096 9318
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 3700 9036 3752 9042
rect 3700 8978 3752 8984
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 848 8968 900 8974
rect 848 8910 900 8916
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 860 8673 888 8910
rect 2964 8900 3016 8906
rect 2964 8842 3016 8848
rect 846 8664 902 8673
rect 846 8599 902 8608
rect 2976 8498 3004 8842
rect 3436 8786 3464 8910
rect 3712 8786 3740 8978
rect 3792 8968 3844 8974
rect 4068 8968 4120 8974
rect 3792 8910 3844 8916
rect 3896 8916 4068 8922
rect 3896 8910 4120 8916
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 3436 8758 3740 8786
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 2700 6866 2728 8434
rect 2780 8356 2832 8362
rect 2780 8298 2832 8304
rect 2792 7410 2820 8298
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2884 7478 2912 7822
rect 2976 7818 3004 8434
rect 3422 8392 3478 8401
rect 3422 8327 3478 8336
rect 2964 7812 3016 7818
rect 2964 7754 3016 7760
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 3436 7206 3464 8327
rect 3528 7954 3556 8758
rect 3804 8634 3832 8910
rect 3896 8894 4108 8910
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3712 8514 3740 8570
rect 3896 8514 3924 8894
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3608 8492 3660 8498
rect 3712 8486 3924 8514
rect 3988 8498 4016 8774
rect 3608 8434 3660 8440
rect 3620 8022 3648 8434
rect 3700 8356 3752 8362
rect 3700 8298 3752 8304
rect 3608 8016 3660 8022
rect 3608 7958 3660 7964
rect 3516 7948 3568 7954
rect 3516 7890 3568 7896
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 1964 6322 1992 6734
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 2148 5302 2176 6802
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2332 6186 2360 6734
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2424 6390 2452 6598
rect 2608 6458 2636 6734
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2412 6384 2464 6390
rect 2412 6326 2464 6332
rect 2872 6384 2924 6390
rect 2872 6326 2924 6332
rect 2320 6180 2372 6186
rect 2320 6122 2372 6128
rect 2884 5778 2912 6326
rect 3068 6322 3096 6666
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 3436 6118 3464 7142
rect 3528 6934 3556 7890
rect 3620 7886 3648 7958
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 3516 6928 3568 6934
rect 3516 6870 3568 6876
rect 3712 6730 3740 8298
rect 3792 8016 3844 8022
rect 3792 7958 3844 7964
rect 3804 6798 3832 7958
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3700 6724 3752 6730
rect 3700 6666 3752 6672
rect 3804 6186 3832 6734
rect 3896 6458 3924 8486
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 4172 8378 4200 8910
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 4080 8350 4200 8378
rect 4264 8362 4292 8434
rect 4448 8401 4476 8434
rect 4434 8392 4490 8401
rect 4252 8356 4304 8362
rect 4080 8090 4108 8350
rect 4434 8327 4490 8336
rect 4252 8298 4304 8304
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 3988 6798 4016 7278
rect 3976 6792 4028 6798
rect 4080 6780 4108 7890
rect 4632 7478 4660 8774
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4896 8560 4948 8566
rect 4896 8502 4948 8508
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4724 8022 4752 8434
rect 4712 8016 4764 8022
rect 4712 7958 4764 7964
rect 4908 7954 4936 8502
rect 5276 8498 5304 8910
rect 5460 8498 5488 8978
rect 5552 8974 5580 9318
rect 7668 9178 7696 10367
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 6932 9081 6960 9114
rect 6918 9072 6974 9081
rect 6918 9007 6974 9016
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 4712 7812 4764 7818
rect 4712 7754 4764 7760
rect 4620 7472 4672 7478
rect 4620 7414 4672 7420
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4436 6792 4488 6798
rect 4080 6752 4436 6780
rect 3976 6734 4028 6740
rect 4436 6734 4488 6740
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 3988 6390 4016 6734
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 3792 6180 3844 6186
rect 3792 6122 3844 6128
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 3436 5710 3464 6054
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 2136 5296 2188 5302
rect 2136 5238 2188 5244
rect 2688 5296 2740 5302
rect 2688 5238 2740 5244
rect 2700 4758 2728 5238
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 2688 4752 2740 4758
rect 2688 4694 2740 4700
rect 2412 4480 2464 4486
rect 2412 4422 2464 4428
rect 2228 4072 2280 4078
rect 2228 4014 2280 4020
rect 2240 3738 2268 4014
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 2240 3602 2268 3674
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 2424 3466 2452 4422
rect 2412 3460 2464 3466
rect 2412 3402 2464 3408
rect 2700 2990 2728 4694
rect 3160 4146 3188 4966
rect 3240 4548 3292 4554
rect 3240 4490 3292 4496
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3252 3058 3280 4490
rect 3344 3194 3372 5170
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 3620 4826 3648 4966
rect 3608 4820 3660 4826
rect 3608 4762 3660 4768
rect 3608 4684 3660 4690
rect 3608 4626 3660 4632
rect 3620 3670 3648 4626
rect 3712 4554 3740 5646
rect 3804 5642 3832 6122
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4724 5914 4752 7754
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 5276 7002 5304 7890
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 5368 6458 5396 8298
rect 5460 7546 5488 8434
rect 5552 8090 5580 8910
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6196 8634 6224 8774
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6656 8498 6684 8774
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 7116 8430 7144 8978
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5644 7342 5672 8230
rect 6196 7478 6224 8230
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 6380 7410 6408 7822
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 6276 7336 6328 7342
rect 6276 7278 6328 7284
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4448 5642 4476 5714
rect 3792 5636 3844 5642
rect 3792 5578 3844 5584
rect 4068 5636 4120 5642
rect 4068 5578 4120 5584
rect 4436 5636 4488 5642
rect 4436 5578 4488 5584
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3988 5166 4016 5510
rect 3976 5160 4028 5166
rect 3896 5108 3976 5114
rect 3896 5102 4028 5108
rect 3896 5086 4016 5102
rect 3896 4826 3924 5086
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 3884 4684 3936 4690
rect 3884 4626 3936 4632
rect 3700 4548 3752 4554
rect 3700 4490 3752 4496
rect 3712 4282 3740 4490
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 3608 3664 3660 3670
rect 3608 3606 3660 3612
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 2688 2984 2740 2990
rect 2688 2926 2740 2932
rect 2700 2378 2728 2926
rect 3252 2514 3280 2994
rect 3240 2508 3292 2514
rect 3240 2450 3292 2456
rect 3344 2446 3372 2994
rect 3620 2990 3648 3606
rect 3700 3460 3752 3466
rect 3700 3402 3752 3408
rect 3608 2984 3660 2990
rect 3608 2926 3660 2932
rect 3712 2582 3740 3402
rect 3700 2576 3752 2582
rect 3700 2518 3752 2524
rect 3332 2440 3384 2446
rect 3332 2382 3384 2388
rect 3804 2378 3832 4422
rect 3896 3738 3924 4626
rect 3988 4622 4016 4966
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 3988 2530 4016 2926
rect 4080 2825 4108 5578
rect 4448 5370 4476 5578
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4528 5296 4580 5302
rect 4580 5256 4660 5284
rect 4528 5238 4580 5244
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4528 4548 4580 4554
rect 4528 4490 4580 4496
rect 4540 3924 4568 4490
rect 4632 4078 4660 5256
rect 4724 4214 4752 5850
rect 4816 5234 4844 6054
rect 4908 5642 4936 6394
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 5000 5710 5028 6258
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5172 6180 5224 6186
rect 5172 6122 5224 6128
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 4896 5636 4948 5642
rect 4896 5578 4948 5584
rect 5184 5574 5212 6122
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 4908 4468 4936 5306
rect 4988 5228 5040 5234
rect 5276 5216 5304 6054
rect 5368 5370 5396 6190
rect 5552 5846 5580 6734
rect 6092 6724 6144 6730
rect 6092 6666 6144 6672
rect 6104 5914 6132 6666
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 6196 5778 6224 7142
rect 6288 5914 6316 7278
rect 6380 6798 6408 7346
rect 7116 6866 7144 8366
rect 7484 7546 7512 8910
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7668 7818 7696 8230
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7838 7712 7894 7721
rect 7838 7647 7894 7656
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7104 6860 7156 6866
rect 7024 6820 7104 6848
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6380 6322 6408 6734
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5040 5188 5304 5216
rect 4988 5170 5040 5176
rect 5000 4554 5028 5170
rect 5080 5092 5132 5098
rect 5080 5034 5132 5040
rect 5264 5092 5316 5098
rect 5264 5034 5316 5040
rect 5092 4826 5120 5034
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 4988 4548 5040 4554
rect 4988 4490 5040 4496
rect 4816 4440 4936 4468
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 4816 4146 4844 4440
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4620 4072 4672 4078
rect 4620 4014 4672 4020
rect 4540 3896 4660 3924
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3720 4660 3896
rect 4804 3732 4856 3738
rect 4632 3692 4804 3720
rect 4804 3674 4856 3680
rect 4344 3392 4396 3398
rect 4344 3334 4396 3340
rect 4356 2990 4384 3334
rect 4816 3040 4844 3674
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4988 3052 5040 3058
rect 4816 3012 4988 3040
rect 4344 2984 4396 2990
rect 4344 2926 4396 2932
rect 4066 2816 4122 2825
rect 4066 2751 4122 2760
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 3988 2502 4200 2530
rect 4816 2514 4844 3012
rect 4988 2994 5040 3000
rect 5276 2582 5304 5034
rect 5368 4826 5396 5306
rect 5552 5166 5580 5646
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5540 4616 5592 4622
rect 5816 4616 5868 4622
rect 5540 4558 5592 4564
rect 5736 4564 5816 4570
rect 5736 4558 5868 4564
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5368 3194 5396 4082
rect 5552 3738 5580 4558
rect 5736 4542 5856 4558
rect 5736 4078 5764 4542
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5736 3942 5764 4014
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 4896 2576 4948 2582
rect 4896 2518 4948 2524
rect 5264 2576 5316 2582
rect 5264 2518 5316 2524
rect 2688 2372 2740 2378
rect 2688 2314 2740 2320
rect 3792 2372 3844 2378
rect 3792 2314 3844 2320
rect 4172 2310 4200 2502
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 4908 2310 4936 2518
rect 5552 2446 5580 3674
rect 5736 3534 5764 3878
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5908 3460 5960 3466
rect 5908 3402 5960 3408
rect 5920 2650 5948 3402
rect 6012 2990 6040 5102
rect 6104 5030 6132 5170
rect 7024 5166 7052 6820
rect 7104 6802 7156 6808
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7116 5778 7144 6598
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7104 5772 7156 5778
rect 7104 5714 7156 5720
rect 7208 5370 7236 6258
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7484 5234 7512 6598
rect 7576 6390 7604 6598
rect 7668 6458 7696 6598
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7564 6384 7616 6390
rect 7564 6326 7616 6332
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 6196 4622 6224 4966
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 7484 3534 7512 4762
rect 7668 4622 7696 6054
rect 7852 5914 7880 7647
rect 7930 6352 7986 6361
rect 7930 6287 7986 6296
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7838 4992 7894 5001
rect 7838 4927 7894 4936
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7748 4548 7800 4554
rect 7748 4490 7800 4496
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 6104 3058 6132 3470
rect 7668 3398 7696 3878
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 5908 2644 5960 2650
rect 5908 2586 5960 2592
rect 6012 2514 6040 2926
rect 6656 2650 6684 2994
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 7116 2514 7144 2790
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7668 2446 7696 3334
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 2964 2304 3016 2310
rect 2964 2246 3016 2252
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 4896 2304 4948 2310
rect 7760 2281 7788 4490
rect 7852 3738 7880 4927
rect 7944 4826 7972 6287
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 7838 3632 7894 3641
rect 7838 3567 7894 3576
rect 7852 2650 7880 3567
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 4896 2246 4948 2252
rect 7746 2272 7802 2281
rect 2976 2106 3004 2246
rect 4874 2204 5182 2213
rect 7746 2207 7802 2216
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 2964 2100 3016 2106
rect 2964 2042 3016 2048
rect 6920 2100 6972 2106
rect 6920 2042 6972 2048
rect 6932 921 6960 2042
rect 6918 912 6974 921
rect 6918 847 6974 856
<< via2 >>
rect 7654 10376 7710 10432
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 846 8608 902 8664
rect 3422 8336 3478 8392
rect 4434 8336 4490 8392
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 6918 9016 6974 9072
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 7838 7656 7894 7712
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4066 2760 4122 2816
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 7930 6296 7986 6352
rect 7838 4936 7894 4992
rect 7838 3576 7894 3632
rect 7746 2216 7802 2272
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 6918 856 6974 912
<< metal3 >>
rect 7649 10434 7715 10437
rect 8595 10434 9395 10464
rect 7649 10432 9395 10434
rect 7649 10376 7654 10432
rect 7710 10376 9395 10432
rect 7649 10374 9395 10376
rect 7649 10371 7715 10374
rect 8595 10344 9395 10374
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 6913 9074 6979 9077
rect 8595 9074 9395 9104
rect 6913 9072 9395 9074
rect 6913 9016 6918 9072
rect 6974 9016 9395 9072
rect 6913 9014 9395 9016
rect 6913 9011 6979 9014
rect 8595 8984 9395 9014
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 841 8666 907 8669
rect 798 8664 907 8666
rect 798 8608 846 8664
rect 902 8608 907 8664
rect 798 8603 907 8608
rect 798 8560 858 8603
rect 0 8470 858 8560
rect 0 8440 800 8470
rect 3417 8394 3483 8397
rect 4429 8394 4495 8397
rect 3417 8392 4495 8394
rect 3417 8336 3422 8392
rect 3478 8336 4434 8392
rect 4490 8336 4495 8392
rect 3417 8334 4495 8336
rect 3417 8331 3483 8334
rect 4429 8331 4495 8334
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 7833 7714 7899 7717
rect 8595 7714 9395 7744
rect 7833 7712 9395 7714
rect 7833 7656 7838 7712
rect 7894 7656 9395 7712
rect 7833 7654 9395 7656
rect 7833 7651 7899 7654
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 8595 7624 9395 7654
rect 4870 7583 5186 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 7925 6354 7991 6357
rect 8595 6354 9395 6384
rect 7925 6352 9395 6354
rect 7925 6296 7930 6352
rect 7986 6296 9395 6352
rect 7925 6294 9395 6296
rect 7925 6291 7991 6294
rect 8595 6264 9395 6294
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 7833 4994 7899 4997
rect 8595 4994 9395 5024
rect 7833 4992 9395 4994
rect 7833 4936 7838 4992
rect 7894 4936 9395 4992
rect 7833 4934 9395 4936
rect 7833 4931 7899 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 8595 4904 9395 4934
rect 4210 4863 4526 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 7833 3634 7899 3637
rect 8595 3634 9395 3664
rect 7833 3632 9395 3634
rect 7833 3576 7838 3632
rect 7894 3576 9395 3632
rect 7833 3574 9395 3576
rect 7833 3571 7899 3574
rect 8595 3544 9395 3574
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 0 2818 800 2848
rect 4061 2818 4127 2821
rect 0 2816 4127 2818
rect 0 2760 4066 2816
rect 4122 2760 4127 2816
rect 0 2758 4127 2760
rect 0 2728 800 2758
rect 4061 2755 4127 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 7741 2274 7807 2277
rect 8595 2274 9395 2304
rect 7741 2272 9395 2274
rect 7741 2216 7746 2272
rect 7802 2216 9395 2272
rect 7741 2214 9395 2216
rect 7741 2211 7807 2214
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 8595 2184 9395 2214
rect 4870 2143 5186 2144
rect 6913 914 6979 917
rect 8595 914 9395 944
rect 6913 912 9395 914
rect 6913 856 6918 912
rect 6974 856 9395 912
rect 6913 854 9395 856
rect 6913 851 6979 854
rect 8595 824 9395 854
<< via3 >>
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 9280 4528 9296
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 8736 5188 9296
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__nand2b_2  _31_
timestamp -3599
transform 1 0 3036 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _32_
timestamp -3599
transform -1 0 2944 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _33_
timestamp -3599
transform 1 0 2668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _34_
timestamp -3599
transform 1 0 3128 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _35_
timestamp -3599
transform 1 0 3864 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _36_
timestamp -3599
transform -1 0 4140 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _37_
timestamp -3599
transform 1 0 3220 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _38_
timestamp -3599
transform 1 0 4876 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _39_
timestamp -3599
transform -1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _40_
timestamp 1562532584
transform -1 0 4416 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _41_
timestamp -3599
transform 1 0 2668 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _42_
timestamp -3599
transform 1 0 1840 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _43_
timestamp -3599
transform 1 0 2392 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _44_
timestamp -3599
transform -1 0 3680 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _45_
timestamp -3599
transform -1 0 4692 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _46_
timestamp -3599
transform -1 0 5612 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _47_
timestamp -3599
transform -1 0 2760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _48_
timestamp -3599
transform -1 0 4692 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _49_
timestamp -3599
transform -1 0 4232 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _50_
timestamp -3599
transform -1 0 4048 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _51_
timestamp -3599
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _52_
timestamp -3599
transform 1 0 4232 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_4  _53_
timestamp -3599
transform -1 0 3772 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_1  _54_
timestamp -3599
transform 1 0 6624 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _55_
timestamp -3599
transform -1 0 5980 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _56_
timestamp -3599
transform 1 0 5428 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _57_
timestamp -3599
transform 1 0 6348 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _58_
timestamp -3599
transform 1 0 7176 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _59_
timestamp -3599
transform -1 0 6256 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _60_
timestamp -3599
transform -1 0 7268 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _61_
timestamp -3599
transform 1 0 6624 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _62_
timestamp -3599
transform 1 0 2208 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _63_
timestamp -3599
transform 1 0 2392 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _64_
timestamp -3599
transform 1 0 3864 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _65_
timestamp -3599
transform 1 0 4140 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _66_
timestamp -3599
transform 1 0 2760 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _67_
timestamp -3599
transform 1 0 2484 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _68_
timestamp -3599
transform 1 0 3864 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _69_
timestamp -3599
transform 1 0 3956 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _70_
timestamp -3599
transform 1 0 6348 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _71_
timestamp -3599
transform 1 0 5980 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _72_
timestamp -3599
transform 1 0 6348 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _73_
timestamp -3599
transform 1 0 6072 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _74_
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _75_
timestamp -3599
transform 1 0 5704 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _76_
timestamp -3599
transform -1 0 8004 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _77_
timestamp -3599
transform 1 0 6348 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _78_
timestamp -3599
transform 1 0 1564 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp -3599
transform 1 0 4048 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp -3599
transform 1 0 4416 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp -3599
transform 1 0 4692 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  clkload0
timestamp -3599
transform 1 0 5336 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3
timestamp -3599
transform 1 0 1380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11
timestamp -3599
transform 1 0 2116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29
timestamp -3599
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -3599
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp -3599
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69
timestamp -3599
transform 1 0 7452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3
timestamp -3599
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_11
timestamp -3599
transform 1 0 2116 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_73
timestamp -3599
transform 1 0 7820 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp -3599
transform 1 0 1380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_11
timestamp -3599
transform 1 0 2116 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp -3599
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_52
timestamp -3599
transform 1 0 5888 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_69
timestamp -3599
transform 1 0 7452 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp -3599
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_11
timestamp -3599
transform 1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_30
timestamp -3599
transform 1 0 3864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_73
timestamp -3599
transform 1 0 7820 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp -3599
transform 1 0 1380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_11
timestamp -3599
transform 1 0 2116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_49
timestamp -3599
transform 1 0 5612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_70
timestamp -3599
transform 1 0 7544 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3
timestamp -3599
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_11
timestamp -3599
transform 1 0 2116 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_5_28
timestamp -3599
transform 1 0 3680 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_47
timestamp -3599
transform 1 0 5428 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_74
timestamp -3599
transform 1 0 7912 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp -3599
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_11
timestamp -3599
transform 1 0 2116 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_19
timestamp -3599
transform 1 0 2852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_29
timestamp -3599
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_52
timestamp -3599
transform 1 0 5888 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_70
timestamp -3599
transform 1 0 7544 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3
timestamp -3599
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_11
timestamp -3599
transform 1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_39
timestamp -3599
transform 1 0 4692 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_73
timestamp -3599
transform 1 0 7820 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7
timestamp -3599
transform 1 0 1748 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp -3599
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_49
timestamp -3599
transform 1 0 5612 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp -3599
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_11
timestamp -3599
transform 1 0 2116 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_73
timestamp -3599
transform 1 0 7820 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp -3599
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_11
timestamp -3599
transform 1 0 2116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_39
timestamp -3599
transform 1 0 4692 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp -3599
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_6
timestamp -3599
transform 1 0 1656 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_14
timestamp -3599
transform 1 0 2392 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_29
timestamp -3599
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_57
timestamp -3599
transform 1 0 6348 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_73
timestamp -3599
transform 1 0 7820 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp -3599
transform 1 0 3220 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp -3599
transform 1 0 3956 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp -3599
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp -3599
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp -3599
transform -1 0 7912 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp -3599
transform 1 0 5520 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp -3599
transform 1 0 7268 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp -3599
transform 1 0 4784 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp -3599
transform 1 0 5520 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp -3599
transform 1 0 3956 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp -3599
transform 1 0 4692 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp -3599
transform -1 0 7544 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp -3599
transform -1 0 6808 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp -3599
transform 1 0 4416 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp -3599
transform -1 0 5520 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp -3599
transform -1 0 3680 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp -3599
transform 1 0 2208 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp -3599
transform -1 0 4692 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp -3599
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp -3599
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output2
timestamp -3599
transform -1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp -3599
transform 1 0 5704 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp -3599
transform 1 0 7636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp -3599
transform 1 0 7636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp -3599
transform 1 0 7636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp -3599
transform 1 0 7636 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp -3599
transform -1 0 3128 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp -3599
transform 1 0 7452 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_13
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_14
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 8280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_15
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 8280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_16
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 8280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_17
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 8280 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_18
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 8280 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_19
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 8280 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_20
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 8280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_21
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 8280 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_22
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 8280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_23
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 8280 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_24
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 8280 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_25
timestamp -3599
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -3599
transform -1 0 8280 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_28
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_29
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_30
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_31
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_32
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_33
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_34
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_35
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_36
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_37
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_38
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_39
timestamp -3599
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_40
timestamp -3599
transform 1 0 6256 0 1 8704
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 9296 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 9296 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 8595 824 9395 944 0 FreeSans 480 0 0 0 counter_out[0]
port 3 nsew signal output
flabel metal3 s 8595 2184 9395 2304 0 FreeSans 480 0 0 0 counter_out[1]
port 4 nsew signal output
flabel metal3 s 8595 3544 9395 3664 0 FreeSans 480 0 0 0 counter_out[2]
port 5 nsew signal output
flabel metal3 s 8595 4904 9395 5024 0 FreeSans 480 0 0 0 counter_out[3]
port 6 nsew signal output
flabel metal3 s 8595 6264 9395 6384 0 FreeSans 480 0 0 0 counter_out[4]
port 7 nsew signal output
flabel metal3 s 8595 7624 9395 7744 0 FreeSans 480 0 0 0 counter_out[5]
port 8 nsew signal output
flabel metal3 s 8595 8984 9395 9104 0 FreeSans 480 0 0 0 counter_out[6]
port 9 nsew signal output
flabel metal3 s 8595 10344 9395 10464 0 FreeSans 480 0 0 0 counter_out[7]
port 10 nsew signal output
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 trigger
port 11 nsew signal input
rlabel metal1 4692 8704 4692 8704 0 VGND
rlabel metal1 4692 9248 4692 9248 0 VPWR
rlabel viali 2525 3502 2525 3502 0 _00_
rlabel metal2 3174 4556 3174 4556 0 _01_
rlabel metal1 3680 2550 3680 2550 0 _02_
rlabel metal1 4222 4590 4222 4590 0 _03_
rlabel metal1 2392 6154 2392 6154 0 _04_
rlabel metal2 2806 7854 2806 7854 0 _05_
rlabel metal1 3940 6698 3940 6698 0 _06_
rlabel metal1 4457 7446 4457 7446 0 _07_
rlabel via1 6665 3026 6665 3026 0 _08_
rlabel metal1 6102 3434 6102 3434 0 _09_
rlabel metal1 4830 2924 4830 2924 0 _10_
rlabel metal1 5658 5100 5658 5100 0 _11_
rlabel metal1 7636 5202 7636 5202 0 _12_
rlabel metal1 6440 5746 6440 5746 0 _13_
rlabel metal1 7314 8364 7314 8364 0 _14_
rlabel metal1 6164 8466 6164 8466 0 _15_
rlabel metal2 2714 2652 2714 2652 0 _16_
rlabel metal1 3174 3162 3174 3162 0 _17_
rlabel metal1 3680 2618 3680 2618 0 _18_
rlabel metal1 3650 2346 3650 2346 0 _19_
rlabel metal1 2898 5066 2898 5066 0 _20_
rlabel metal2 1978 6528 1978 6528 0 _21_
rlabel metal1 4462 4046 4462 4046 0 _22_
rlabel metal2 2438 6494 2438 6494 0 _23_
rlabel metal1 4600 5814 4600 5814 0 _24_
rlabel metal1 2530 8500 2530 8500 0 _25_
rlabel metal2 2714 7650 2714 7650 0 _26_
rlabel via1 3818 8942 3818 8942 0 _27_
rlabel metal2 4002 8636 4002 8636 0 _28_
rlabel metal1 4462 8908 4462 8908 0 _29_
rlabel metal2 5658 7786 5658 7786 0 _30_
rlabel metal2 4094 4199 4094 4199 0 clk
rlabel metal1 5060 5882 5060 5882 0 clknet_0_clk
rlabel metal1 2346 4046 2346 4046 0 clknet_1_0__leaf_clk
rlabel metal1 2530 7412 2530 7412 0 clknet_1_1__leaf_clk
rlabel metal1 6302 2550 6302 2550 0 counter\[0\]
rlabel metal1 3818 4522 3818 4522 0 counter\[1\]
rlabel metal1 5060 3706 5060 3706 0 counter\[2\]
rlabel metal1 5198 5338 5198 5338 0 counter\[3\]
rlabel metal1 6118 6358 6118 6358 0 counter\[4\]
rlabel metal1 3956 6086 3956 6086 0 counter\[5\]
rlabel metal1 4830 8534 4830 8534 0 counter\[6\]
rlabel metal2 5474 8738 5474 8738 0 counter\[7\]
rlabel metal2 2990 2176 2990 2176 0 counter_out[0]
rlabel metal3 8242 2244 8242 2244 0 counter_out[1]
rlabel metal3 8288 3604 8288 3604 0 counter_out[2]
rlabel metal2 7866 4335 7866 4335 0 counter_out[3]
rlabel metal1 7912 4794 7912 4794 0 counter_out[4]
rlabel metal2 7866 6783 7866 6783 0 counter_out[5]
rlabel metal1 4922 9146 4922 9146 0 counter_out[6]
rlabel metal2 7682 9775 7682 9775 0 counter_out[7]
rlabel metal1 2185 8806 2185 8806 0 net1
rlabel metal1 5520 2822 5520 2822 0 net10
rlabel metal1 6486 5202 6486 5202 0 net11
rlabel metal1 6292 4590 6292 4590 0 net12
rlabel metal1 6946 6426 6946 6426 0 net13
rlabel metal2 7222 5814 7222 5814 0 net14
rlabel metal1 6486 8602 6486 8602 0 net15
rlabel via1 7686 7786 7686 7786 0 net16
rlabel metal1 6302 8874 6302 8874 0 net17
rlabel metal1 6424 7446 6424 7446 0 net18
rlabel metal1 5290 3094 5290 3094 0 net19
rlabel metal1 3266 2414 3266 2414 0 net2
rlabel metal2 5382 3638 5382 3638 0 net20
rlabel metal1 6578 5882 6578 5882 0 net21
rlabel metal2 6118 6290 6118 6290 0 net22
rlabel metal1 5290 2278 5290 2278 0 net23
rlabel metal1 4738 9044 4738 9044 0 net24
rlabel metal2 2622 6596 2622 6596 0 net25
rlabel via1 3077 6290 3077 6290 0 net26
rlabel metal1 4048 8058 4048 8058 0 net27
rlabel metal2 3634 4896 3634 4896 0 net28
rlabel metal1 5060 2414 5060 2414 0 net3
rlabel metal1 6026 3366 6026 3366 0 net4
rlabel metal1 6808 4794 6808 4794 0 net5
rlabel metal1 6716 6086 6716 6086 0 net6
rlabel metal1 7268 5746 7268 5746 0 net7
rlabel metal2 5566 9146 5566 9146 0 net8
rlabel metal1 7498 9010 7498 9010 0 net9
rlabel metal3 751 8500 751 8500 0 trigger
rlabel metal2 3634 8160 3634 8160 0 trigger_prev
<< properties >>
string FIXED_BBOX 0 0 9395 11539
<< end >>
