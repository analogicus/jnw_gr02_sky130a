magic
tech sky130A
timestamp 1744492486
<< locali >>
rect -4458 1175 2272 1178
rect -4458 1085 -4261 1175
rect -4171 1085 -2061 1175
rect -1971 1085 1539 1175
rect 1629 1085 2272 1175
rect -4458 1082 2272 1085
rect -4456 1002 -4360 1082
rect -3624 1002 -3528 1082
rect -1424 988 -1328 1082
rect -1056 982 -960 1082
rect -224 964 -128 1082
rect 144 972 240 1082
rect 976 992 1072 1082
rect 1344 992 1440 1082
rect 2176 988 2272 1082
rect -2256 -1292 -2160 -1060
rect -1424 -1292 -1328 -1042
rect -1056 -1292 -960 -1060
rect -224 -1292 -128 -1060
rect 144 -1292 240 -1060
rect 976 -1292 1072 -1060
rect 1344 -1292 1440 -1060
rect 2176 -1292 2272 -1060
rect -2160 -1295 2272 -1292
rect -2160 -1382 -2061 -1295
rect -2256 -1385 -2061 -1382
rect -1971 -1385 -861 -1295
rect -771 -1385 339 -1295
rect 429 -1385 1539 -1295
rect 1629 -1385 2272 -1295
rect -2256 -1388 2272 -1385
rect -2256 -1636 -2160 -1388
rect -4538 -1692 -2160 -1636
rect -2256 -1698 -2160 -1692
<< viali >>
rect -4261 1085 -4171 1175
rect -2061 1085 -1971 1175
rect 1539 1085 1629 1175
rect -4345 -225 -4255 -135
rect -4134 -240 -4020 -120
rect -3587 -237 -3473 -123
rect -3378 -240 -3258 -126
rect -2877 -237 -2763 -123
rect -2617 -237 -2503 -123
rect -2256 -1382 -2160 -1292
rect -2061 -1385 -1971 -1295
rect -861 -1385 -771 -1295
rect 339 -1385 429 -1295
rect 1539 -1385 1629 -1295
<< metal1 >>
rect -3816 1232 432 1328
rect -4264 1175 -4168 1181
rect -4264 1085 -4261 1175
rect -4171 1085 -4168 1175
rect -4264 912 -4168 1085
rect -3816 948 -3720 1232
rect -2064 1175 -1968 1181
rect -2064 1085 -2061 1175
rect -1971 1085 -1968 1175
rect -4328 584 -4296 716
rect -4326 566 -4294 569
rect -4326 531 -4294 534
rect -4264 512 -4168 778
rect -3769 534 -3766 565
rect -3734 534 -3731 565
rect -3818 208 -3722 338
rect -4348 112 -3722 208
rect -4348 -135 -4252 112
rect -3730 -60 -2760 60
rect -4348 -225 -4345 -135
rect -4255 -225 -4252 -135
rect -4348 -231 -4252 -225
rect -4137 -120 -4017 -114
rect -3730 -120 -3610 -60
rect -4137 -240 -4134 -120
rect -4020 -123 -3467 -120
rect -2880 -123 -2760 -60
rect -4020 -237 -3587 -123
rect -3473 -237 -3467 -123
rect -4020 -240 -3467 -237
rect -3384 -126 -3252 -123
rect -3384 -240 -3378 -126
rect -3258 -240 -3252 -126
rect -4137 -246 -4017 -240
rect -3384 -243 -3252 -240
rect -2880 -237 -2877 -123
rect -2763 -237 -2760 -123
rect -2880 -243 -2760 -237
rect -2620 -123 -2500 -117
rect -2620 -237 -2617 -123
rect -2503 -237 -2500 -123
rect -3378 -300 -3258 -243
rect -2620 -300 -2500 -237
rect -2128 -246 -2096 776
rect -3378 -420 -2500 -300
rect -2064 -358 -1968 1085
rect -1616 -268 -1520 848
rect -864 832 -768 1232
rect 336 872 432 1232
rect 1536 1175 1632 1181
rect 1536 1085 1539 1175
rect 1629 1085 1632 1175
rect 1536 892 1632 1085
rect -928 276 -896 766
rect -1226 244 -896 276
rect -928 -206 -896 244
rect -864 -218 -768 748
rect -416 -238 -320 848
rect 272 276 304 746
rect -16 244 304 276
rect 272 -216 304 244
rect -2620 -1270 -2500 -420
rect -2128 -614 -2096 -484
rect -1616 -584 -1520 -402
rect -1616 -614 -1586 -584
rect -2128 -616 -1586 -614
rect -1554 -616 -1520 -584
rect -2128 -646 -1520 -616
rect -416 -634 -320 -412
rect 336 -438 432 828
rect -1616 -918 -1520 -646
rect -928 -666 -320 -634
rect 784 -644 880 828
rect 1472 -246 1504 756
rect 1536 -448 1632 818
rect 1194 -584 1226 -581
rect 1472 -584 1504 -484
rect 1226 -616 1504 -584
rect 1984 -592 2080 828
rect 1194 -619 1226 -616
rect -928 -788 -896 -666
rect -416 -878 -320 -666
rect 272 -676 1504 -644
rect 272 -788 304 -676
rect 784 -898 880 -676
rect 1472 -788 1504 -676
rect 1984 -688 2468 -592
rect 1984 -908 2080 -688
rect -2128 -1174 -2096 -1084
rect -2128 -1209 -2096 -1206
rect -2620 -1289 -2160 -1270
rect -2620 -1292 -2154 -1289
rect -2620 -1382 -2256 -1292
rect -2160 -1382 -2154 -1292
rect -2620 -1385 -2154 -1382
rect -2064 -1295 -1968 -984
rect -928 -1134 -896 -1084
rect -928 -1174 -894 -1134
rect -929 -1206 -926 -1174
rect -894 -1206 -891 -1174
rect -2064 -1385 -2061 -1295
rect -1971 -1385 -1968 -1295
rect -2620 -1390 -2160 -1385
rect -2064 -1391 -1968 -1385
rect -864 -1295 -768 -984
rect -864 -1385 -861 -1295
rect -771 -1385 -768 -1295
rect -864 -1391 -768 -1385
rect 336 -1295 432 -984
rect 336 -1385 339 -1295
rect 429 -1385 432 -1295
rect 336 -1391 432 -1385
rect 1536 -1295 1632 -984
rect 1536 -1385 1539 -1295
rect 1629 -1385 1632 -1295
rect 1536 -1391 1632 -1385
<< via1 >>
rect -4326 534 -4294 566
rect -3766 534 -3734 565
rect -1586 -616 -1554 -584
rect 1194 -616 1226 -584
rect -2128 -1206 -2096 -1174
rect -926 -1206 -894 -1174
<< metal2 >>
rect -3766 566 -3734 568
rect -4329 534 -4326 566
rect -4294 565 -3734 566
rect -4294 534 -3766 565
rect -3766 531 -3734 534
rect -1589 -616 -1586 -584
rect -1554 -616 1194 -584
rect 1226 -616 1229 -584
rect -926 -1174 -894 -1171
rect -2131 -1206 -2128 -1174
rect -2096 -1206 -926 -1174
rect -926 -1209 -894 -1206
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_0 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 -1008 0 1 -536
box -92 -64 924 464
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_1
timestamp 1740610800
transform 1 0 192 0 1 664
box -92 -64 924 464
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_2
timestamp 1740610800
transform 1 0 -1008 0 1 -136
box -92 -64 924 464
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_3
timestamp 1740610800
transform 1 0 -1008 0 1 664
box -92 -64 924 464
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_4
timestamp 1740610800
transform 1 0 -1008 0 1 264
box -92 -64 924 464
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_5
timestamp 1740610800
transform 1 0 192 0 1 -536
box -92 -64 924 464
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_6
timestamp 1740610800
transform 1 0 192 0 1 -136
box -92 -64 924 464
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_7
timestamp 1740610800
transform 1 0 192 0 1 264
box -92 -64 924 464
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_0 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 1392 0 1 -536
box -92 -64 924 464
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_1
timestamp 1740610800
transform 1 0 -2208 0 -1 264
box -92 -64 924 464
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_2
timestamp 1740610800
transform 1 0 -2208 0 1 -536
box -92 -64 924 464
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_3
timestamp 1740610800
transform 1 0 -2208 0 1 264
box -92 -64 924 464
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_4
timestamp 1740610800
transform 1 0 -2208 0 1 664
box -92 -64 924 464
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_5
timestamp 1740610800
transform 1 0 1392 0 1 664
box -92 -64 924 464
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_6
timestamp 1740610800
transform 1 0 1392 0 1 -136
box -92 -64 924 464
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_7
timestamp 1740610800
transform 1 0 1392 0 1 264
box -92 -64 924 464
use JNWTR_RPPO2  JNWTR_RPPO2_0 ../JNW_TR_SKY130A
timestamp 1744284492
transform -1 0 -3076 0 1 -1700
box 0 0 724 1720
use JNWTR_RPPO2  JNWTR_RPPO2_1
timestamp 1744284492
transform -1 0 -2316 0 1 -1700
box 0 0 724 1720
use JNWTR_RPPO2  x6
timestamp 1744284492
transform -1 0 -3836 0 1 -1700
box 0 0 724 1720
use JNWATR_PCH_12C5F0  xa01
timestamp 1740610800
transform 1 0 -4408 0 1 264
box -92 -64 924 464
use JNWATR_PCH_12C5F0  xa02
timestamp 1740610800
transform 1 0 -4408 0 1 664
box -92 -64 924 464
use JNWATR_NCH_12C5F0  xc01 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 -1008 0 1 -1136
box -92 -64 924 464
use JNWATR_NCH_12C5F0  xc02
timestamp 1740610800
transform 1 0 -2208 0 1 -1136
box -92 -64 924 464
use JNWATR_NCH_12C5F0  xc03
timestamp 1740610800
transform 1 0 1392 0 1 -1136
box -92 -64 924 464
use JNWATR_NCH_12C5F0  xc04
timestamp 1740610800
transform 1 0 192 0 1 -1136
box -92 -64 924 464
<< labels >>
flabel metal1 -1226 244 -1194 276 0 FreeSans 800 0 0 0 VIP
port 6 nsew
flabel metal1 -16 244 16 276 0 FreeSans 800 0 0 0 VIN
port 7 nsew
flabel locali -1424 -1388 -1328 -1292 0 FreeSans 800 0 0 0 VSS
port 8 nsew
flabel locali -2828 1082 -2732 1178 0 FreeSans 800 0 0 0 VDD
port 11 nsew
flabel metal1 2372 -688 2468 -592 0 FreeSans 800 0 0 0 VOUT
port 12 nsew
<< properties >>
string FIXED_BBOX 0 0 1172 3620
<< end >>
