*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/JNW_CURRENT_lpe.spi
#else
.include ../../../work/xsch/JNW_CURRENT.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3 method=gear

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD VSS dc 1.8 


*V4 V_M4P VSS dc 0.5
V5 V_M5P VSS dc 0.5

*V6 V_BIAS VSS dc 0.7
*V7 V_REF VSS dc 1.2

*R1P V_M1P V_M1N 1m

*R2P V_M2P V_M2N 1m

*R3P V_M3P V_M3N 1m

*R4P V_M4P VSS 1m

*R5P V_M5P VSS 1m

R6P V_BIAS VSS 1MEG

*R7P V_REF VSS 1MEG

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all 


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

*optran 0 0 0 1n 1u 0


tran 1n 100n 1n
write
quit


.endc

.end
