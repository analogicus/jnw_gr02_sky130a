*Automatic generated instance fron ../../tech/scripts/genxdut dig
adut [clk
+ n_rst
+ trigger
+ ]
+ [reset
+ counter_out.7
+ counter_out.6
+ counter_out.5
+ counter_out.4
+ counter_out.3
+ counter_out.2
+ counter_out.1
+ counter_out.0
+ counter.7
+ counter.6
+ counter.5
+ counter.4
+ counter.3
+ counter.2
+ counter.1
+ counter.0
+ ] null dut
.model dut d_cosim simulation="../dig.so" delay=10p queue_size=8096

* Inputs
Rsvi0 clk 0 1G
Rsvi1 n_rst 0 1G
Rsvi2 trigger 0 1G

* Outputs
Rsvi3 reset 0 1G
Rsvi4 counter_out.7 0 1G
Rsvi5 counter_out.6 0 1G
Rsvi6 counter_out.5 0 1G
Rsvi7 counter_out.4 0 1G
Rsvi8 counter_out.3 0 1G
Rsvi9 counter_out.2 0 1G
Rsvi10 counter_out.1 0 1G
Rsvi11 counter_out.0 0 1G
Rsvi12 counter.7 0 1G
Rsvi13 counter.6 0 1G
Rsvi14 counter.5 0 1G
Rsvi15 counter.4 0 1G
Rsvi16 counter.3 0 1G
Rsvi17 counter.2 0 1G
Rsvi18 counter.1 0 1G
Rsvi19 counter.0 0 1G

.save v(reset)

E_STATE_counter_out dec_counter_out 0 value={( 0 
+ + 128*v(counter_out.7)/AVDD
+ + 64*v(counter_out.6)/AVDD
+ + 32*v(counter_out.5)/AVDD
+ + 16*v(counter_out.4)/AVDD
+ + 8*v(counter_out.3)/AVDD
+ + 4*v(counter_out.2)/AVDD
+ + 2*v(counter_out.1)/AVDD
+ + 1*v(counter_out.0)/AVDD
+)/1000}
.save v(dec_counter_out)

E_STATE_counter dec_counter 0 value={( 0 
+ + 128*v(counter.7)/AVDD
+ + 64*v(counter.6)/AVDD
+ + 32*v(counter.5)/AVDD
+ + 16*v(counter.4)/AVDD
+ + 8*v(counter.3)/AVDD
+ + 4*v(counter.2)/AVDD
+ + 2*v(counter.1)/AVDD
+ + 1*v(counter.0)/AVDD
+)/1000}
.save v(dec_counter)

