*Automatic generated instance fron ../../tech/scripts/genxdut dig
adut [clk
+ trigger
+ ]
+ [counter_out.7
+ counter_out.6
+ counter_out.5
+ counter_out.4
+ counter_out.3
+ counter_out.2
+ counter_out.1
+ counter_out.0
+ ] null dut
.model dut d_cosim simulation="../dig.so" delay=10p queue_size=8096

* Inputs
Rsvi0 clk 0 1G
Rsvi1 trigger 0 1G

* Outputs
Rsvi2 counter_out.7 0 1G
Rsvi3 counter_out.6 0 1G
Rsvi4 counter_out.5 0 1G
Rsvi5 counter_out.4 0 1G
Rsvi6 counter_out.3 0 1G
Rsvi7 counter_out.2 0 1G
Rsvi8 counter_out.1 0 1G
Rsvi9 counter_out.0 0 1G

E_STATE_counter_out dec_counter_out 0 value={( 0 
+ + 128*v(counter_out.7)/AVDD
+ + 64*v(counter_out.6)/AVDD
+ + 32*v(counter_out.5)/AVDD
+ + 16*v(counter_out.4)/AVDD
+ + 8*v(counter_out.3)/AVDD
+ + 4*v(counter_out.2)/AVDD
+ + 2*v(counter_out.1)/AVDD
+ + 1*v(counter_out.0)/AVDD
+)/1000}
.save v(dec_counter_out)

