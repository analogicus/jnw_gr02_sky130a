magic
tech sky130A
magscale 1 2
timestamp 1745878851
<< locali >>
rect -9716 2350 4544 2356
rect -9716 2170 -9322 2350
rect -9142 2170 -4122 2350
rect -3942 2170 3078 2350
rect 3258 2170 4544 2350
rect -9716 2164 4544 2170
rect -9712 2004 -9520 2164
rect -8048 2004 -7856 2164
rect -2848 1976 -2656 2164
rect -2112 1964 -1920 2164
rect -448 1928 -256 2164
rect 288 1944 480 2164
rect 1952 1984 2144 2164
rect 2688 1984 2880 2164
rect 4352 1976 4544 2164
rect -4512 -2584 -4320 -2120
rect -2848 -2584 -2656 -2084
rect -2112 -2584 -1920 -2120
rect -448 -2584 -256 -2120
rect 288 -2584 480 -2120
rect 1952 -2584 2144 -2120
rect 2688 -2584 2880 -2120
rect 4352 -2584 4544 -2120
rect -4516 -2590 4544 -2584
rect -4516 -2770 -4122 -2590
rect -3942 -2770 -1722 -2590
rect -1542 -2770 678 -2590
rect 858 -2770 3078 -2590
rect 3258 -2770 4544 -2590
rect -4516 -2776 4544 -2770
rect -4512 -3204 -4320 -2776
rect -9796 -3396 -4320 -3204
<< viali >>
rect -9322 2170 -9142 2350
rect -4122 2170 -3942 2350
rect 3078 2170 3258 2350
rect -9430 -470 -9250 -290
rect -8956 -480 -8716 -240
rect -7634 -474 -7406 -246
rect -7156 -480 -6916 -240
rect -5974 -474 -5746 -246
rect -5414 -474 -5186 -246
rect -4122 -2770 -3942 -2590
rect -1722 -2770 -1542 -2590
rect 678 -2770 858 -2590
rect 3078 -2770 3258 -2590
<< metal1 >>
rect -8432 2464 864 2656
rect -9328 2350 -9136 2362
rect -9328 2170 -9322 2350
rect -9142 2170 -9136 2350
rect -9456 1138 -9392 1824
rect -9456 1132 -9388 1138
rect -9456 1068 -9452 1132
rect -9456 1062 -9388 1068
rect -9456 864 -9392 1062
rect -9328 736 -9136 2170
rect -8432 1376 -8240 2464
rect -4128 2350 -3936 2362
rect -4128 2170 -4122 2350
rect -3942 2170 -3936 2350
rect -8432 376 -8240 896
rect -9436 184 -8240 376
rect -9436 -290 -9244 184
rect -7874 40 -5740 280
rect -9436 -470 -9430 -290
rect -9250 -470 -9244 -290
rect -9436 -482 -9244 -470
rect -8987 -240 -8468 -232
rect -7874 -240 -7634 40
rect -7188 -240 -6667 -231
rect -8987 -480 -8956 -240
rect -8716 -246 -7380 -240
rect -8716 -474 -7634 -246
rect -7406 -474 -7380 -246
rect -8716 -480 -7380 -474
rect -7188 -480 -7156 -240
rect -6916 -480 -6300 -240
rect -8987 -487 -8468 -480
rect -7188 -488 -6667 -480
rect -6540 -580 -6300 -480
rect -5980 -246 -5740 40
rect -5980 -474 -5974 -246
rect -5746 -474 -5740 -246
rect -5980 -486 -5740 -474
rect -5420 -246 -5180 -234
rect -5420 -474 -5414 -246
rect -5186 -474 -5180 -246
rect -5420 -580 -5180 -474
rect -6540 -820 -5180 -580
rect -5420 -2520 -5180 -820
rect -4256 -1228 -4192 1552
rect -4128 -716 -3936 2170
rect -3232 -1168 -3040 1696
rect -1856 552 -1792 1824
rect -2452 488 -1792 552
rect -1856 -992 -1792 488
rect -1728 -992 -1536 2464
rect -3232 -1228 -3172 -1168
rect -4256 -1232 -3172 -1228
rect -3108 -1232 -3040 -1168
rect -4256 -1292 -3040 -1232
rect -832 -1268 -640 1824
rect 544 552 608 1952
rect -32 488 608 552
rect 544 -864 608 488
rect 672 -876 864 2464
rect 3072 2350 3264 2362
rect 3072 2170 3078 2350
rect 3258 2170 3264 2350
rect -3232 -1836 -3040 -1292
rect -1856 -1332 -640 -1268
rect 1568 -1288 1760 2016
rect 2388 -1168 2452 -1162
rect 2944 -1168 3008 1888
rect 3072 -896 3264 2170
rect 2452 -1232 3008 -1168
rect 3968 -1184 4160 1888
rect 2388 -1238 2452 -1232
rect -4256 -2348 -4192 -1952
rect -4256 -2418 -4192 -2412
rect -4128 -2520 -3936 -1968
rect -1856 -2268 -1792 -1332
rect -832 -1756 -640 -1332
rect 544 -1352 3008 -1288
rect 544 -1760 608 -1352
rect 1568 -1796 1760 -1352
rect 2944 -1760 3008 -1352
rect 3968 -1376 4936 -1184
rect -1856 -2348 -1788 -2268
rect -1858 -2412 -1852 -2348
rect -1788 -2412 -1782 -2348
rect -5420 -2590 -3936 -2520
rect -5420 -2760 -4122 -2590
rect -4128 -2770 -4122 -2760
rect -3942 -2770 -3936 -2590
rect -4128 -2782 -3936 -2770
rect -1728 -2590 -1536 -1968
rect -1728 -2770 -1722 -2590
rect -1542 -2770 -1536 -2590
rect -1728 -2782 -1536 -2770
rect 672 -2590 864 -1968
rect 672 -2770 678 -2590
rect 858 -2770 864 -2590
rect 672 -2782 864 -2770
rect 3072 -2590 3264 -1568
rect 3968 -2144 4160 -1376
rect 3072 -2770 3078 -2590
rect 3258 -2770 3264 -2590
rect 3072 -2782 3264 -2770
<< via1 >>
rect -9452 1068 -9388 1132
rect -8332 1068 -8268 1130
rect -3172 -1232 -3108 -1168
rect 2388 -1232 2452 -1168
rect -4256 -2412 -4192 -2348
rect -1852 -2412 -1788 -2348
<< metal2 >>
rect -8332 1132 -8268 1136
rect -9458 1068 -9452 1132
rect -9388 1130 -8268 1132
rect -9388 1068 -8332 1130
rect -8332 1062 -8268 1068
rect -3178 -1232 -3172 -1168
rect -3108 -1232 2388 -1168
rect 2452 -1232 2458 -1168
rect -1852 -2348 -1788 -2342
rect -4262 -2412 -4256 -2348
rect -4192 -2412 -1852 -2348
rect -1852 -2418 -1788 -2412
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_0 ../JNW_ATR_SKY130A
timestamp 1745878851
transform 1 0 -2016 0 1 -1072
box -184 -128 1848 928
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_1
timestamp 1745878851
transform 1 0 384 0 1 1328
box -184 -128 1848 928
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_2
timestamp 1745878851
transform 1 0 -2016 0 1 -272
box -184 -128 1848 928
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_3
timestamp 1745878851
transform 1 0 -2016 0 1 1328
box -184 -128 1848 928
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_4
timestamp 1745878851
transform 1 0 -2016 0 1 528
box -184 -128 1848 928
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_5
timestamp 1745878851
transform 1 0 384 0 1 -1072
box -184 -128 1848 928
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_6
timestamp 1745878851
transform 1 0 384 0 1 -272
box -184 -128 1848 928
use JNWATR_PCH_12C1F2  JNWATR_PCH_12C1F2_7
timestamp 1745878851
transform 1 0 384 0 1 528
box -184 -128 1848 928
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_0 ../JNW_ATR_SKY130A
timestamp 1745878851
transform 1 0 2784 0 1 -1072
box -184 -128 1848 928
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_1
timestamp 1745878851
transform 1 0 -4416 0 -1 528
box -184 -128 1848 928
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_2
timestamp 1745878851
transform 1 0 -4416 0 1 -1072
box -184 -128 1848 928
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_3
timestamp 1745878851
transform 1 0 -4416 0 1 528
box -184 -128 1848 928
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_4
timestamp 1745878851
transform 1 0 -4416 0 1 1328
box -184 -128 1848 928
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_5
timestamp 1745878851
transform 1 0 2784 0 1 1328
box -184 -128 1848 928
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_6
timestamp 1745878851
transform 1 0 2784 0 1 -272
box -184 -128 1848 928
use JNWATR_PCH_12C5F0  JNWATR_PCH_12C5F0_7
timestamp 1745878851
transform 1 0 2784 0 1 528
box -184 -128 1848 928
use JNWTR_RPPO2  JNWTR_RPPO2_0 ../JNW_TR_SKY130A
timestamp 1745878851
transform -1 0 -8352 0 1 -3400
box 0 0 1448 3440
use JNWTR_RPPO2  JNWTR_RPPO2_1
timestamp 1745878851
transform -1 0 -4832 0 1 -3400
box 0 0 1448 3440
use JNWTR_RPPO2  JNWTR_RPPO2_2
timestamp 1745878851
transform -1 0 -6552 0 1 -3400
box 0 0 1448 3440
use JNWATR_PCH_12C5F0  xa01
timestamp 1745878851
transform 1 0 -9616 0 1 528
box -184 -128 1848 928
use JNWATR_PCH_12C5F0  xa02
timestamp 1745878851
transform 1 0 -9616 0 1 1328
box -184 -128 1848 928
use JNWATR_NCH_12C5F0  xc01 ../JNW_ATR_SKY130A
timestamp 1745878851
transform 1 0 -2016 0 1 -2272
box -184 -128 1848 928
use JNWATR_NCH_12C5F0  xc02
timestamp 1745878851
transform 1 0 -4416 0 1 -2272
box -184 -128 1848 928
use JNWATR_NCH_12C5F0  xc03
timestamp 1745878851
transform 1 0 2784 0 1 -2272
box -184 -128 1848 928
use JNWATR_NCH_12C5F0  xc04
timestamp 1745878851
transform 1 0 384 0 1 -2272
box -184 -128 1848 928
<< labels >>
flabel metal1 -2452 488 -2388 552 0 FreeSans 1600 0 0 0 VIP
port 6 nsew
flabel metal1 -32 488 32 552 0 FreeSans 1600 0 0 0 VIN
port 7 nsew
flabel locali -2848 -2776 -2656 -2584 0 FreeSans 1600 0 0 0 VSS
port 8 nsew
flabel locali -5656 2164 -5464 2356 0 FreeSans 1600 0 0 0 VDD
port 11 nsew
flabel metal1 4744 -1376 4936 -1184 0 FreeSans 1600 0 0 0 VOUT
port 12 nsew
<< properties >>
string FIXED_BBOX 0 0 2344 7240
<< end >>
