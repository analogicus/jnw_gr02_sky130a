VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dig
  CLASS BLOCK ;
  FOREIGN dig ;
  ORIGIN 0.000 0.000 ;
  SIZE 33.000 BY 120.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 109.040 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 109.040 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 0.300 29.200 ;
    END
  END clk
  PIN counter_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 32.700 6.840 33.000 7.440 ;
    END
  END counter_out[0]
  PIN counter_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 32.700 21.800 33.000 22.400 ;
    END
  END counter_out[1]
  PIN counter_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 32.700 36.760 33.000 37.360 ;
    END
  END counter_out[2]
  PIN counter_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 32.700 51.720 33.000 52.320 ;
    END
  END counter_out[3]
  PIN counter_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 32.700 66.680 33.000 67.280 ;
    END
  END counter_out[4]
  PIN counter_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 32.700 81.640 33.000 82.240 ;
    END
  END counter_out[5]
  PIN counter_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 32.700 96.600 33.000 97.200 ;
    END
  END counter_out[6]
  PIN counter_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 32.700 111.560 33.000 112.160 ;
    END
  END counter_out[7]
  PIN trigger
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 0.300 89.040 ;
    END
  END trigger
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 27.330 108.885 ;
      LAYER li1 ;
        RECT 5.520 10.795 27.140 108.885 ;
      LAYER met1 ;
        RECT 3.290 10.640 32.130 109.040 ;
      LAYER met2 ;
        RECT 3.310 6.955 32.110 112.045 ;
      LAYER met3 ;
        RECT 0.300 111.160 32.300 112.025 ;
        RECT 0.300 97.600 32.700 111.160 ;
        RECT 0.300 96.200 32.300 97.600 ;
        RECT 0.300 89.440 32.700 96.200 ;
        RECT 0.700 88.040 32.700 89.440 ;
        RECT 0.300 82.640 32.700 88.040 ;
        RECT 0.300 81.240 32.300 82.640 ;
        RECT 0.300 67.680 32.700 81.240 ;
        RECT 0.300 66.280 32.300 67.680 ;
        RECT 0.300 52.720 32.700 66.280 ;
        RECT 0.300 51.320 32.300 52.720 ;
        RECT 0.300 37.760 32.700 51.320 ;
        RECT 0.300 36.360 32.300 37.760 ;
        RECT 0.300 29.600 32.700 36.360 ;
        RECT 0.700 28.200 32.700 29.600 ;
        RECT 0.300 22.800 32.700 28.200 ;
        RECT 0.300 21.400 32.300 22.800 ;
        RECT 0.300 7.840 32.700 21.400 ;
        RECT 0.300 6.975 32.300 7.840 ;
  END
END dig
END LIBRARY

