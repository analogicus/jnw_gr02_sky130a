magic
tech sky130A
magscale 1 2
timestamp 1744566493
<< locali >>
rect 23804 -1010 33016 -1004
rect 23804 -1190 25078 -1010
rect 25258 -1190 33016 -1010
rect 23804 -1196 33016 -1190
rect 24688 -2224 24880 -1196
rect 26352 -2224 26544 -1196
rect 32120 -1458 32296 -1196
rect 27820 -1550 29170 -1490
rect 24688 -7250 24880 -4920
rect 26352 -5304 26544 -4872
rect 26096 -5496 26556 -5304
rect 26096 -5672 26288 -5496
rect 24688 -7430 24690 -7250
rect 24870 -7430 24880 -7250
rect 24688 -8644 24880 -7430
rect 26096 -8644 26288 -6884
rect 22220 -8836 26288 -8644
rect 24688 -10024 24880 -8836
rect 26840 -9260 27060 -1970
rect 27820 -2610 27880 -1550
rect 27280 -3130 27340 -2790
rect 28540 -3130 28600 -2810
rect 27280 -3142 28600 -3130
rect 27280 -3190 28540 -3142
rect 27820 -3970 27880 -3190
rect 27280 -4530 27340 -4230
rect 28540 -4530 28600 -4230
rect 27280 -4542 28600 -4530
rect 27280 -4590 28540 -4542
rect 27820 -5450 27880 -4590
rect 27280 -5970 27340 -5610
rect 28540 -5970 28600 -5630
rect 27280 -5982 28600 -5970
rect 27280 -6030 28540 -5982
rect 27820 -6870 27880 -6030
rect 27280 -7370 27340 -7030
rect 28540 -7370 28600 -7030
rect 27280 -7382 28600 -7370
rect 27280 -7430 28540 -7382
rect 27820 -8270 27880 -7430
rect 27280 -8770 27340 -8410
rect 28540 -8770 28600 -8410
rect 28840 -8720 29020 -1838
rect 29110 -5430 29170 -1550
rect 32120 -1622 32126 -1458
rect 32290 -1622 32296 -1458
rect 32120 -1628 32296 -1622
rect 31670 -2010 31880 -1950
rect 30844 -4898 31036 -2164
rect 31820 -2630 31880 -2010
rect 31280 -3250 31340 -2830
rect 32540 -3250 32600 -2810
rect 31280 -3310 32600 -3250
rect 31820 -3970 31880 -3310
rect 31280 -4490 31340 -4150
rect 32540 -4490 32600 -4170
rect 32824 -4436 33016 -1196
rect 31280 -4496 32600 -4490
rect 31280 -4544 31956 -4496
rect 32004 -4544 32600 -4496
rect 31280 -4550 32600 -4544
rect 30844 -5062 30858 -4898
rect 31022 -5062 31036 -4898
rect 29110 -5490 29862 -5430
rect 29110 -8770 29170 -5490
rect 27280 -8782 29170 -8770
rect 27280 -8830 28540 -8782
rect 28600 -8830 29170 -8782
rect 26840 -9390 27060 -9380
rect 30844 -10024 31036 -5062
rect 24688 -10216 31036 -10024
<< viali >>
rect 25078 -1190 25258 -1010
rect 24690 -7430 24870 -7250
rect 28840 -1838 29020 -1670
rect 28540 -3190 28600 -3142
rect 28540 -4590 28600 -4542
rect 28540 -6030 28600 -5982
rect 28540 -7430 28600 -7382
rect 32126 -1622 32290 -1458
rect 31956 -4544 32004 -4496
rect 30858 -5062 31022 -4898
rect 29862 -5490 29910 -5430
rect 28540 -8830 28600 -8782
rect 26840 -9380 27060 -9260
<< metal1 >>
rect 25072 -1010 25264 -998
rect 25072 -1190 25078 -1010
rect 25258 -1190 25264 -1010
rect 25072 -2356 25264 -1190
rect 32120 -1458 32296 -1446
rect 32120 -1622 32126 -1458
rect 32290 -1622 32296 -1458
rect 25968 -1670 29036 -1664
rect 25968 -1672 28840 -1670
rect 25968 -1848 28120 -1672
rect 28296 -1838 28840 -1672
rect 29020 -1838 29036 -1670
rect 32120 -1692 32296 -1622
rect 28296 -1848 29036 -1838
rect 25968 -1856 29036 -1848
rect 25968 -2316 26160 -1856
rect 32114 -1868 32120 -1692
rect 32296 -1868 32302 -1692
rect 24944 -3092 25008 -2708
rect 25072 -3176 25264 -2408
rect 28528 -3142 28612 -3136
rect 28528 -3190 28540 -3142
rect 28600 -3190 28612 -3142
rect 28528 -3196 28612 -3190
rect 28540 -3230 28600 -3196
rect 28540 -3296 28600 -3290
rect 24944 -3768 25008 -3468
rect 25968 -3640 26160 -3424
rect 25968 -3768 26496 -3640
rect 24944 -3832 26496 -3768
rect 24364 -4236 26156 -4044
rect 24364 -4312 24556 -4236
rect 23624 -4504 24556 -4312
rect 24944 -4412 25008 -4236
rect 25964 -4496 26156 -4236
rect 24944 -6412 25008 -4968
rect 25072 -7244 25264 -4608
rect 26304 -5304 26496 -3832
rect 31950 -4496 32010 -4484
rect 28528 -4542 28612 -4536
rect 28528 -4590 28540 -4542
rect 28600 -4590 28612 -4542
rect 28528 -4596 28612 -4590
rect 31950 -4544 31956 -4496
rect 32004 -4544 32010 -4496
rect 28540 -4630 28600 -4596
rect 28540 -4696 28600 -4690
rect 31352 -4892 31528 -4886
rect 30846 -4898 31352 -4892
rect 30846 -5062 30858 -4898
rect 31022 -5062 31352 -4898
rect 30846 -5068 31352 -5062
rect 31352 -5074 31528 -5068
rect 25712 -5496 26496 -5304
rect 29856 -5430 29916 -5418
rect 31950 -5430 32010 -4544
rect 29856 -5490 29862 -5430
rect 29910 -5490 32010 -5430
rect 25712 -5704 25904 -5496
rect 29856 -5502 29916 -5490
rect 28528 -5982 28612 -5976
rect 28528 -6030 28540 -5982
rect 28600 -6030 28612 -5982
rect 28528 -6036 28612 -6030
rect 28540 -6070 28600 -6036
rect 28540 -6136 28600 -6130
rect 24678 -7250 25264 -7244
rect 24678 -7430 24690 -7250
rect 24870 -7430 25264 -7250
rect 24678 -7436 25264 -7430
rect 22888 -8092 23012 -8028
rect 22888 -8412 22952 -8092
rect 25712 -9245 25904 -6444
rect 28528 -7382 28612 -7376
rect 28528 -7430 28540 -7382
rect 28600 -7430 28612 -7382
rect 28528 -7436 28612 -7430
rect 28540 -7470 28600 -7436
rect 28540 -7536 28600 -7530
rect 28528 -8782 28612 -8776
rect 28528 -8830 28540 -8782
rect 28600 -8830 28612 -8782
rect 28528 -8836 28612 -8830
rect 28540 -8870 28600 -8836
rect 28540 -8936 28600 -8930
rect 25712 -9260 27285 -9245
rect 25712 -9376 26840 -9260
rect 25725 -9380 26840 -9376
rect 27060 -9380 27285 -9260
rect 25725 -9395 27285 -9380
rect 27435 -9395 27441 -9245
rect 20892 -15784 21084 -14744
rect 20684 -15976 21084 -15784
<< via1 >>
rect 28120 -1848 28296 -1672
rect 32120 -1868 32296 -1692
rect 28540 -3290 28600 -3230
rect 28540 -4690 28600 -4630
rect 31352 -5068 31528 -4892
rect 28540 -6130 28600 -6070
rect 28540 -7530 28600 -7470
rect 28540 -8930 28600 -8870
rect 27285 -9395 27435 -9245
<< metal2 >>
rect 28120 -1672 28296 -1666
rect 28120 -1957 28296 -1848
rect 32120 -1692 32296 -1686
rect 32120 -1937 32296 -1868
rect 28116 -2123 28125 -1957
rect 28291 -2123 28300 -1957
rect 32116 -2103 32125 -1937
rect 32291 -2103 32300 -1937
rect 32120 -2108 32296 -2103
rect 28120 -2128 28296 -2123
rect 28534 -3290 28540 -3230
rect 28600 -3290 28606 -3230
rect 28540 -3330 28600 -3290
rect 28381 -3390 28390 -3330
rect 28446 -3390 28600 -3330
rect 28534 -4690 28540 -4630
rect 28600 -4690 28606 -4630
rect 28540 -4730 28600 -4690
rect 28381 -4790 28390 -4730
rect 28446 -4790 28600 -4730
rect 31585 -4892 31751 -4888
rect 31346 -5068 31352 -4892
rect 31528 -4897 31756 -4892
rect 31528 -5063 31585 -4897
rect 31751 -5063 31756 -4897
rect 31528 -5068 31756 -5063
rect 31585 -5072 31751 -5068
rect 28534 -6130 28540 -6070
rect 28600 -6130 28606 -6070
rect 28540 -6170 28600 -6130
rect 28381 -6230 28390 -6170
rect 28446 -6230 28600 -6170
rect 28534 -7530 28540 -7470
rect 28600 -7530 28606 -7470
rect 28540 -7570 28600 -7530
rect 28381 -7630 28390 -7570
rect 28446 -7630 28600 -7570
rect 28534 -8930 28540 -8870
rect 28600 -8930 28606 -8870
rect 28540 -8970 28600 -8930
rect 28381 -9030 28390 -8970
rect 28446 -9030 28600 -8970
rect 27285 -9245 27435 -9239
rect 27435 -9395 27615 -9245
rect 27755 -9395 27764 -9245
rect 27285 -9401 27435 -9395
<< via2 >>
rect 28125 -2123 28291 -1957
rect 32125 -2103 32291 -1937
rect 28390 -3390 28446 -3330
rect 28390 -4790 28446 -4730
rect 31585 -5063 31751 -4897
rect 28390 -6230 28446 -6170
rect 28390 -7630 28446 -7570
rect 28390 -9030 28446 -8970
rect 27615 -9395 27755 -9245
<< metal3 >>
rect 32120 -1937 32296 -1932
rect 28120 -1957 28296 -1952
rect 28120 -2123 28125 -1957
rect 28291 -2123 28296 -1957
rect 27580 -9240 27756 -2692
rect 28120 -8652 28296 -2123
rect 32120 -2103 32125 -1937
rect 32291 -2103 32296 -1937
rect 28385 -3330 28451 -3325
rect 28385 -3390 28390 -3330
rect 28446 -3390 29750 -3330
rect 28385 -3395 28451 -3390
rect 28385 -4730 28451 -4725
rect 28385 -4790 28390 -4730
rect 28446 -4790 29770 -4730
rect 28385 -4795 28451 -4790
rect 31580 -4897 31756 -2852
rect 32120 -3888 32296 -2103
rect 31580 -5063 31585 -4897
rect 31751 -5063 31756 -4897
rect 31580 -5068 31756 -5063
rect 28385 -6170 28451 -6165
rect 28385 -6230 28390 -6170
rect 28446 -6230 29870 -6170
rect 28385 -6235 28451 -6230
rect 28385 -7570 28451 -7565
rect 28385 -7630 28390 -7570
rect 28446 -7630 29830 -7570
rect 28385 -7635 28451 -7630
rect 28385 -8970 28451 -8965
rect 28385 -9030 28390 -8970
rect 28446 -9030 29890 -8970
rect 28385 -9035 28451 -9030
rect 27580 -9245 27760 -9240
rect 27580 -9395 27615 -9245
rect 27755 -9395 27847 -9245
rect 27995 -9395 28001 -9245
rect 27580 -9400 27760 -9395
rect 27580 -9408 27756 -9400
<< via3 >>
rect 27847 -9395 27995 -9245
<< metal4 >>
rect 27846 -9245 27996 -9244
rect 30185 -9245 30335 -3695
rect 27846 -9395 27847 -9245
rect 27995 -9395 30335 -9245
rect 27846 -9396 27996 -9395
use JNWTR_CAPX1  JNWTR_CAPX1_0 ../JNW_TR_SKY130A
timestamp 1737500400
transform 0 1 29500 1 0 -9720
box 0 0 1080 1080
use JNWTR_IVX4_CV  JNWTR_IVX4_CV_0 ../JNW_TR_SKY130A
timestamp 1744538702
transform 1 0 26950 0 1 -8680
box -150 -120 2130 920
use JNWTR_IVX4_CV  JNWTR_IVX4_CV_1
timestamp 1744538702
transform 1 0 26950 0 1 -4380
box -150 -120 2130 920
use JNWTR_IVX4_CV  JNWTR_IVX4_CV_2
timestamp 1744538702
transform 1 0 26950 0 1 -7180
box -150 -120 2130 920
use JNWTR_IVX4_CV  JNWTR_IVX4_CV_3
timestamp 1744538702
transform 1 0 26950 0 1 -5880
box -150 -120 2130 920
use JNWTR_IVX4_CV  JNWTR_IVX4_CV_4
timestamp 1744538702
transform 1 0 26950 0 1 -2980
box -150 -120 2130 920
use JNW_VIS_TI  x2 ../JNW_GR02_SKY130A
timestamp 1744548984
transform 1 0 14388 0 1 1400
box -9344 -19400 9900 -2398
use JNWTR_CAPX1  x7
timestamp 1737500400
transform 0 -1 30580 1 0 -3800
box 0 0 1080 1080
use JNWATR_NCH_8C1F2  x8 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 24784 0 1 -7072
box -184 -128 1592 928
use JNWATR_NCH_12C1F2  x9 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 24784 0 1 -5072
box -184 -128 1848 928
use JNWTR_IVX4_CV  x10
timestamp 1744538702
transform 1 0 30950 0 1 -3080
box -150 -120 2130 920
use JNWATR_NCH_8C1F2  x11
timestamp 1734044400
transform 1 0 24784 0 1 -6272
box -184 -128 1592 928
use JNWATR_PCH_12C1F2  x12 ../JNW_ATR_SKY130A
timestamp 1744535236
transform 1 0 24784 0 1 -3672
box -184 -128 1848 928
use JNWATR_PCH_12C1F2  x13
timestamp 1744535236
transform 1 0 24784 0 1 -2872
box -184 -128 1848 928
use JNWTR_IVX4_CV  x14
timestamp 1744538702
transform 1 0 30950 0 1 -4420
box -150 -120 2130 920
use JNWTR_CAPX1  x15
timestamp 1737500400
transform 0 -1 30580 1 0 -5300
box 0 0 1080 1080
use JNWTR_CAPX1  x16
timestamp 1737500400
transform 0 -1 30580 1 0 -6800
box 0 0 1080 1080
use JNWTR_CAPX1  x17
timestamp 1737500400
transform 0 -1 30580 1 0 -8300
box 0 0 1080 1080
<< labels >>
flabel locali 24688 -10216 31036 -10024 0 FreeSans 1600 0 0 0 VSS
port 0 nsew
flabel locali 31670 -2010 31730 -1950 0 FreeSans 1600 0 0 0 VOUT
port 1 nsew
flabel metal1 22948 -8092 23012 -8028 0 FreeSans 1600 0 0 0 PWR_UP
port 2 nsew
flabel locali 27324 -1196 27516 -1004 0 FreeSans 1600 0 0 0 VDD
port 3 nsew
flabel space 7184 -7156 7376 -6964 0 FreeSans 1600 0 0 0 VREF
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 34124 12080
<< end >>
