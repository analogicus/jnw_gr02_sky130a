** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_GR02_SKY130A/TB_JNW_VIS_ITIME.sch
**.subckt TB_JNW_VIS_ITIME VDD VSS PWR_UP RST VOUT LPI LPO ITEMP_O ITEMP_I
*.ipin VDD
*.ipin VSS
*.ipin PWR_UP
*.ipin RST
*.opin VOUT
*.opin LPI
*.opin LPO
*.opin ITEMP_O
*.ipin ITEMP_I
x1 VDD VREF VOUT ITEMP_I RST VSS JNW_VIS_ITIME
x2 VDD VREF LPI LPO ITEMP_O PWR_UP VSS JNW_VIS_TI
**.ends

* expanding   symbol:  JNW_GR02_SKY130A/JNW_VIS_ITIME.sym # of pins=6
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_GR02_SKY130A/JNW_VIS_ITIME.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_GR02_SKY130A/JNW_VIS_ITIME.sch
.subckt JNW_VIS_ITIME VDD VREF VOUT I_TEMP RST VSS
*.ipin VDD
*.ipin VSS
*.ipin VREF
*.ipin I_TEMP
*.ipin RST
*.opin VOUT
x7 VDD I_TEMP VREF VSS VOUT JNW_VIS_OTA
x4 I_TEMP RST VSS VSS JNWATR_NCH_8C1F2
x1<0> I_TEMP VSS JNWTR_CAPX1
x1<1> I_TEMP VSS JNWTR_CAPX1
x1<2> I_TEMP VSS JNWTR_CAPX1
x1<3> I_TEMP VSS JNWTR_CAPX1
x1<4> I_TEMP VSS JNWTR_CAPX1
x1<5> I_TEMP VSS JNWTR_CAPX1
x1<6> I_TEMP VSS JNWTR_CAPX1
x1<7> I_TEMP VSS JNWTR_CAPX1
x1<8> I_TEMP VSS JNWTR_CAPX1
x1<9> I_TEMP VSS JNWTR_CAPX1
x1<10> I_TEMP VSS JNWTR_CAPX1
x1<11> I_TEMP VSS JNWTR_CAPX1
x1<12> I_TEMP VSS JNWTR_CAPX1
x1<13> I_TEMP VSS JNWTR_CAPX1
x1<14> I_TEMP VSS JNWTR_CAPX1
x1<15> I_TEMP VSS JNWTR_CAPX1
x1<16> I_TEMP VSS JNWTR_CAPX1
x1<17> I_TEMP VSS JNWTR_CAPX1
x1<18> I_TEMP VSS JNWTR_CAPX1
x1<19> I_TEMP VSS JNWTR_CAPX1
x1<20> I_TEMP VSS JNWTR_CAPX1
x1<21> I_TEMP VSS JNWTR_CAPX1
x1<22> I_TEMP VSS JNWTR_CAPX1
x1<23> I_TEMP VSS JNWTR_CAPX1
x1<24> I_TEMP VSS JNWTR_CAPX1
x1<25> I_TEMP VSS JNWTR_CAPX1
x1<26> I_TEMP VSS JNWTR_CAPX1
x1<27> I_TEMP VSS JNWTR_CAPX1
x1<28> I_TEMP VSS JNWTR_CAPX1
x1<29> I_TEMP VSS JNWTR_CAPX1
x1<30> I_TEMP VSS JNWTR_CAPX1
x1<31> I_TEMP VSS JNWTR_CAPX1
x1<32> I_TEMP VSS JNWTR_CAPX1
x1<33> I_TEMP VSS JNWTR_CAPX1
x1<34> I_TEMP VSS JNWTR_CAPX1
x1<35> I_TEMP VSS JNWTR_CAPX1
x1<36> I_TEMP VSS JNWTR_CAPX1
x1<37> I_TEMP VSS JNWTR_CAPX1
x1<38> I_TEMP VSS JNWTR_CAPX1
x1<39> I_TEMP VSS JNWTR_CAPX1
x1<40> I_TEMP VSS JNWTR_CAPX1
x1<41> I_TEMP VSS JNWTR_CAPX1
x1<42> I_TEMP VSS JNWTR_CAPX1
x1<43> I_TEMP VSS JNWTR_CAPX1
x1<44> I_TEMP VSS JNWTR_CAPX1
x1<45> I_TEMP VSS JNWTR_CAPX1
x1<46> I_TEMP VSS JNWTR_CAPX1
x1<47> I_TEMP VSS JNWTR_CAPX1
x1<48> I_TEMP VSS JNWTR_CAPX1
x1<49> I_TEMP VSS JNWTR_CAPX1
x1<50> I_TEMP VSS JNWTR_CAPX1
x1<51> I_TEMP VSS JNWTR_CAPX1
x1<52> I_TEMP VSS JNWTR_CAPX1
x1<53> I_TEMP VSS JNWTR_CAPX1
x1<54> I_TEMP VSS JNWTR_CAPX1
x1<55> I_TEMP VSS JNWTR_CAPX1
x1<56> I_TEMP VSS JNWTR_CAPX1
x1<57> I_TEMP VSS JNWTR_CAPX1
x1<58> I_TEMP VSS JNWTR_CAPX1
x1<59> I_TEMP VSS JNWTR_CAPX1
x1<60> I_TEMP VSS JNWTR_CAPX1
x1<61> I_TEMP VSS JNWTR_CAPX1
x1<62> I_TEMP VSS JNWTR_CAPX1
x1<63> I_TEMP VSS JNWTR_CAPX1
x1<64> I_TEMP VSS JNWTR_CAPX1
x1<65> I_TEMP VSS JNWTR_CAPX1
x1<66> I_TEMP VSS JNWTR_CAPX1
x1<67> I_TEMP VSS JNWTR_CAPX1
x1<68> I_TEMP VSS JNWTR_CAPX1
x1<69> I_TEMP VSS JNWTR_CAPX1
x1<70> I_TEMP VSS JNWTR_CAPX1
x1<71> I_TEMP VSS JNWTR_CAPX1
x1<72> I_TEMP VSS JNWTR_CAPX1
x1<73> I_TEMP VSS JNWTR_CAPX1
x1<74> I_TEMP VSS JNWTR_CAPX1
x1<75> I_TEMP VSS JNWTR_CAPX1
x1<76> I_TEMP VSS JNWTR_CAPX1
x1<77> I_TEMP VSS JNWTR_CAPX1
x1<78> I_TEMP VSS JNWTR_CAPX1
x1<79> I_TEMP VSS JNWTR_CAPX1
x1<80> I_TEMP VSS JNWTR_CAPX1
x1<81> I_TEMP VSS JNWTR_CAPX1
x1<82> I_TEMP VSS JNWTR_CAPX1
x1<83> I_TEMP VSS JNWTR_CAPX1
x1<84> I_TEMP VSS JNWTR_CAPX1
x1<85> I_TEMP VSS JNWTR_CAPX1
x1<86> I_TEMP VSS JNWTR_CAPX1
x1<87> I_TEMP VSS JNWTR_CAPX1
x1<88> I_TEMP VSS JNWTR_CAPX1
x1<89> I_TEMP VSS JNWTR_CAPX1
x1<90> I_TEMP VSS JNWTR_CAPX1
x1<91> I_TEMP VSS JNWTR_CAPX1
x1<92> I_TEMP VSS JNWTR_CAPX1
x1<93> I_TEMP VSS JNWTR_CAPX1
x1<94> I_TEMP VSS JNWTR_CAPX1
x1<95> I_TEMP VSS JNWTR_CAPX1
x1<96> I_TEMP VSS JNWTR_CAPX1
x1<97> I_TEMP VSS JNWTR_CAPX1
x1<98> I_TEMP VSS JNWTR_CAPX1
x1<99> I_TEMP VSS JNWTR_CAPX1
.ends


* expanding   symbol:  JNW_GR02_SKY130A/JNW_VIS_TI.sym # of pins=7
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_GR02_SKY130A/JNW_VIS_TI.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_GR02_SKY130A/JNW_VIS_TI.sch
.subckt JNW_VIS_TI VDD VREF LPI LPO I_TEMP PWR_UP VSS
*.ipin VDD
*.ipin VSS
*.opin VREF
*.opin I_TEMP
*.ipin PWR_UP
*.opin LPI
*.opin LPO
XQ1 VSS VSS VIN sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1 mult=1
XQ2 VSS VSS VD2 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=8 mult=8
x7 VDD VIN VIP VSS LPO JNW_VIS_OTA
x11 VDD PWR_UP LPI VSS JNWATR_NCH_2C1F2
x1<0> LPI VSS JNWTR_CAPX1
x1<1> LPI VSS JNWTR_CAPX1
x1<2> LPI VSS JNWTR_CAPX1
x5<0> VIP VREF VSS JNWTR_RPPO16
x8<0> VD2 VIP VSS JNWTR_RPPO4
x8<1> VD2 VIP VSS JNWTR_RPPO4
x2<0> net1 net1 VDD VDD JNWATR_PCH_8C5F0
x2<1> net1 net1 VDD VDD JNWATR_PCH_8C5F0
x3<0> VIN net1 VDD VDD JNWATR_PCH_8C5F0
x3<1> VIN net1 VDD VDD JNWATR_PCH_8C5F0
x4<0> VREF net1 VDD VDD JNWATR_PCH_8C5F0
x4<1> VREF net1 VDD VDD JNWATR_PCH_8C5F0
x4 I_TEMP net1 VDD VDD JNWATR_PCH_8C5F0
x6 net1 LPI VSS VSS JNWATR_NCH_2C5F0
.ends


* expanding   symbol:  JNW_GR02_SKY130A/JNW_VIS_OTA.sym # of pins=5
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_GR02_SKY130A/JNW_VIS_OTA.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_GR02_SKY130A/JNW_VIS_OTA.sch
.subckt JNW_VIS_OTA VDD VIN VIP VSS VOUT
*.ipin VDD
*.ipin VIP
*.ipin VIN
*.ipin VSS
*.opin VOUT
x1 V2 VIP VOP VOP JNWATR_PCH_2C1F2
x10 V1 VIN VOP VOP JNWATR_PCH_2C1F2
x3 VOUT V1 VSS VSS JNWATR_NCH_2C5F0
x4 V2 V2 VSS VSS JNWATR_NCH_4C5F0
x5 net1 V2 VSS VSS JNWATR_NCH_2C5F0
x6 V1 V1 VSS VSS JNWATR_NCH_4C5F0
x7 VOUT net1 VDD VDD JNWATR_PCH_8C5F0
x8<0> VOP VGS_M VDD VDD JNWATR_PCH_4C1F2
x8<1> VOP VGS_M VDD VDD JNWATR_PCH_4C1F2
x9 VGS_M VGS_M VDD VDD JNWATR_PCH_4C1F2
x11 net1 net1 VDD VDD JNWATR_PCH_8C5F0
x2<0> VSS net2 VSS JNWTR_RPPO8
x1<0> net2 VGS_M VSS JNWTR_RPPO16
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_8C1F2.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_8C1F2.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_8C1F2.sch
.subckt JNWATR_NCH_8C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.22 W=5.76 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_CAPX1.sym # of pins=2
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sch
.subckt JNWTR_CAPX1 A B
*.iopin A
*.iopin B
XC1 B A sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_2C1F2.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_2C1F2.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_2C1F2.sch
.subckt JNWATR_NCH_2C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.22 W=1.92 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RPPO16.sym # of pins=3
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO16.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO16.sch
.subckt JNWTR_RPPO16 N P B
*.iopin P
*.iopin N
*.iopin B
XXA1 N P B JNWTR_RES16
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RPPO4.sym # of pins=3
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO4.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO4.sch
.subckt JNWTR_RPPO4 N P B
*.iopin P
*.iopin N
*.iopin B
XXA1 N P B JNWTR_RES4
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_8C5F0.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_8C5F0.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_8C5F0.sch
.subckt JNWATR_PCH_8C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.94 W=5.76 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_2C5F0.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_2C5F0.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_2C5F0.sch
.subckt JNWATR_NCH_2C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.94 W=1.92 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_2C1F2.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_2C1F2.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_2C1F2.sch
.subckt JNWATR_PCH_2C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.22 W=1.92 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sch
.subckt JNWATR_NCH_4C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.94 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_4C1F2.sym # of pins=4
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C1F2.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C1F2.sch
.subckt JNWATR_PCH_4C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.22 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RPPO8.sym # of pins=3
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO8.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO8.sch
.subckt JNWTR_RPPO8 N P B
*.iopin P
*.iopin N
*.iopin B
XXA1 N P B JNWTR_RES8
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RES16.sym # of pins=3
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RES16.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RES16.sch
.subckt JNWTR_RES16 N P B
*.iopin N
*.iopin P
*.iopin B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_1 INT_1 INT_0 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_2 INT_2 INT_1 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_3 INT_3 INT_2 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_4 INT_4 INT_3 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_5 INT_5 INT_4 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_6 INT_6 INT_5 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_7 INT_7 INT_6 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_8 INT_8 INT_7 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_9 INT_9 INT_8 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_10 INT_10 INT_9 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_11 INT_11 INT_10 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_12 INT_12 INT_11 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_13 INT_13 INT_12 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_14 INT_14 INT_13 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_15 P INT_14 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RES4.sym # of pins=3
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RES4.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RES4.sch
.subckt JNWTR_RES4 N P B
*.iopin N
*.iopin P
*.iopin B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_1 INT_1 INT_0 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_2 INT_2 INT_1 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_3 P INT_2 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RES8.sym # of pins=3
** sym_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RES8.sym
** sch_path: /home/domen/pro/aicex/ip/jnw_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RES8.sch
.subckt JNWTR_RES8 N P B
*.iopin N
*.iopin P
*.iopin B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_1 INT_1 INT_0 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_2 INT_2 INT_1 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_3 INT_3 INT_2 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_4 INT_4 INT_3 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_5 INT_5 INT_4 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_6 INT_6 INT_5 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_7 P INT_6 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
.ends

.end
