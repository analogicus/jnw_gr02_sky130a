*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/JNW_VIS_TI_lpe.spi
#else
.include ../../../work/xsch/JNW_VIS_TI.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3 method=gear

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD VSS dc 1.8 
VPUP PWR_UP VSS PULSE ( 0 1.8 10NS 1PS 1PS 10NS 1S 1)
VSENS I_TEMP 0 dc 0.5

RSH LPO LPI 1u

.ic V(LPI)=0.5

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all i(VSENS) v(VREF)


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=6
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0

set fend = .raw
#ifdef Nosweep
    option temp=27
    tran 10n 1000n 1p
    write
#else
    foreach vtemp {temp_sweep}
        option temp=$vtemp
        tran 10n 1000n 1p
        write {cicname}_$vtemp$fend
    end
#endif

quit


.endc

.end
