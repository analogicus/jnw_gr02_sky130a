magic
tech sky130A
magscale 1 2
timestamp 1744568593
<< locali >>
rect -4982 11670 -4214 11688
rect -4982 11114 -4950 11670
rect -4394 11114 -4214 11670
rect -4982 10408 -4214 11114
rect 16292 11670 16860 11676
rect 16292 11114 16298 11670
rect 16854 11114 16860 11670
rect 16292 10084 16860 11114
rect 16292 10024 16856 10084
rect 10096 5152 10288 5293
rect 10096 5120 10464 5152
rect 9856 4928 10496 5120
rect 9856 4480 9984 4928
rect 10432 4480 10496 4928
rect 9856 4416 10496 4480
rect 15616 4416 17408 4544
rect 14840 4144 14900 4258
rect 15616 4160 15680 4416
rect 17344 4096 17408 4416
rect 18082 4170 18142 4898
rect 14840 4066 14900 4084
rect 14840 4064 14848 4066
rect 17439 3867 17633 3873
rect 17439 3812 17508 3867
rect 17563 3812 17633 3867
rect 14940 3805 15139 3811
rect 14940 3746 14946 3805
rect 15005 3746 15139 3805
rect 14940 3740 15139 3746
rect 17439 3743 17633 3812
rect 14653 3389 14788 3587
rect 15074 3444 15134 3614
rect 17086 3453 17221 3651
rect 17506 3490 17566 3650
rect 14653 3266 14659 3389
rect 14782 3266 14788 3389
rect 17086 3330 17092 3453
rect 17215 3330 17221 3453
rect 17086 3324 17221 3330
rect 14653 3260 14788 3266
rect -8221 -6953 -7651 -5155
rect -8221 -7511 -8215 -6953
rect -7657 -7511 -7651 -6953
rect -8221 -7517 -7651 -7511
<< viali >>
rect -4950 11114 -4394 11670
rect 16298 11114 16854 11670
rect 9984 4480 10432 4928
rect 18082 4898 18142 4958
rect 14840 4258 14900 4318
rect 16584 4166 16701 4283
rect 17508 3812 17563 3867
rect 14946 3746 15005 3805
rect 14659 3266 14782 3389
rect 17092 3330 17215 3453
rect -8215 -7511 -7657 -6953
<< metal1 >>
rect -4962 11748 -4956 12316
rect -4388 11748 -4382 12316
rect 16286 11748 16292 12316
rect 16860 11748 16866 12316
rect -4956 11670 -4388 11748
rect -4956 11114 -4950 11670
rect -4394 11114 -4388 11670
rect -4956 11102 -4388 11114
rect 16292 11670 16860 11748
rect 16292 11114 16298 11670
rect 16854 11114 16860 11670
rect 16292 11102 16860 11114
rect -14100 4892 -1456 5084
rect 3732 3232 3924 5744
rect 18076 4958 18148 4970
rect 9972 4928 10444 4934
rect 9972 4480 9984 4928
rect 10432 4480 10444 4928
rect 18076 4898 18082 4958
rect 18142 4898 18210 4958
rect 18270 4898 18276 4958
rect 18076 4886 18148 4898
rect 19264 4800 19392 6720
rect 9972 4474 10444 4480
rect 14807 4673 19392 4800
rect 9984 4448 10432 4474
rect 14807 4318 14934 4673
rect 14976 4672 19392 4673
rect 16570 4480 16576 4609
rect 16709 4480 16715 4609
rect 14807 4289 14840 4318
rect 14828 4258 14840 4289
rect 14900 4289 14934 4318
rect 14900 4258 14912 4289
rect 14828 4252 14912 4258
rect 16578 4283 16707 4480
rect 16578 4166 16584 4283
rect 16701 4166 16707 4283
rect 16578 4154 16707 4166
rect 9984 3994 10432 4000
rect 17374 3873 17443 3874
rect 17502 3873 17569 3879
rect 17374 3867 17569 3873
rect 17374 3812 17508 3867
rect 17563 3812 17569 3867
rect 14877 3805 15017 3811
rect 14877 3746 14946 3805
rect 15005 3746 15017 3805
rect 14877 3740 15017 3746
rect 17374 3806 17569 3812
rect 10817 3455 10944 3461
rect 10944 3328 11647 3455
rect 14653 3389 14788 3401
rect 10817 3322 10944 3328
rect 14653 3266 14659 3389
rect 14782 3266 14788 3389
rect 3732 3040 12000 3232
rect 14653 3140 14788 3266
rect 14647 3005 14653 3140
rect 14788 3005 14794 3140
rect 14877 2950 14948 3740
rect 17086 3453 17221 3465
rect 17086 3330 17092 3453
rect 17215 3330 17221 3453
rect 17086 3140 17221 3330
rect 17078 3005 17084 3140
rect 17223 3005 17229 3140
rect 17374 2950 17443 3806
rect 17502 3800 17569 3806
rect 10817 2944 10944 2950
rect 14852 2830 18668 2950
rect 10817 2811 10944 2817
rect 992 -3736 1184 -2912
rect 800 -3928 1184 -3736
rect -8221 -6953 -7651 -6941
rect -8221 -7511 -8215 -6953
rect -7657 -7511 -7651 -6953
rect -8221 -7779 -7651 -7511
rect -8227 -8349 -8221 -7779
rect -7651 -8349 -7645 -7779
rect -15740 -10812 -13892 -10692
rect -14012 -12228 -13892 -10812
rect 18548 -12228 18668 2830
rect -14012 -12348 18668 -12228
rect 18548 -12406 18668 -12348
<< via1 >>
rect -4956 11748 -4388 12316
rect 16292 11748 16860 12316
rect 18210 4898 18270 4958
rect 9984 4000 10432 4448
rect 16576 4480 16709 4609
rect 10817 3328 10944 3455
rect 14653 3005 14788 3140
rect 17084 3005 17223 3140
rect 10817 2817 10944 2944
rect -8221 -8349 -7651 -7779
<< metal2 >>
rect -4956 13017 -4388 13022
rect -4960 12395 -4951 13017
rect -4393 12395 -4384 13017
rect 16292 13015 16860 13020
rect -4956 12316 -4388 12395
rect 16288 12393 16297 13015
rect 16855 12393 16864 13015
rect -4956 11742 -4388 11748
rect 16292 12316 16860 12393
rect 16292 11742 16860 11748
rect 13441 4958 20146 4992
rect 13441 4898 18210 4958
rect 18270 4898 20146 4958
rect 13441 4865 20146 4898
rect 9978 4000 9984 4448
rect 10432 4000 10438 4448
rect 9984 3936 10432 4000
rect -15168 544 -3488 608
rect -15168 448 -15040 544
rect -3552 288 -3488 544
rect 2784 288 2848 3700
rect 9975 3488 9984 3936
rect 10432 3488 10441 3936
rect 10811 3328 10817 3455
rect 10944 3328 10950 3455
rect 10817 2944 10944 3328
rect 13441 2944 13568 4865
rect 19501 4627 19620 4636
rect 16576 4609 16709 4615
rect 18367 4609 18500 4618
rect 15863 4480 15872 4609
rect 16001 4480 16576 4609
rect 16709 4480 18367 4609
rect 18500 4480 19501 4609
rect 16576 4474 16709 4480
rect 18367 4471 18500 4480
rect 19620 4480 19625 4609
rect 19501 4452 19620 4461
rect 19117 3155 19242 3164
rect 14653 3140 14788 3146
rect 15356 3140 15492 3149
rect 17084 3140 17223 3146
rect 17853 3140 17989 3149
rect 14788 3005 15356 3140
rect 15492 3005 17084 3140
rect 17223 3005 17853 3140
rect 17989 3005 19117 3140
rect 14653 2999 14788 3005
rect 15356 2996 15492 3005
rect 17084 2999 17223 3005
rect 17853 2996 17989 3005
rect 19242 3005 19247 3140
rect 19117 2980 19242 2989
rect 10811 2817 10817 2944
rect 10944 2817 13568 2944
rect -3552 224 2848 288
rect -8221 -7779 -7651 -7773
rect -8221 -8744 -7651 -8349
rect -8225 -9304 -8216 -8744
rect -7656 -9304 -7647 -8744
rect -8221 -9309 -7651 -9304
<< via2 >>
rect -4951 12395 -4393 13017
rect 16297 12393 16855 13015
rect 9984 3488 10432 3936
rect 15872 4480 16001 4609
rect 18367 4480 18500 4609
rect 19501 4461 19620 4627
rect 15356 3005 15492 3140
rect 17853 3005 17989 3140
rect 19117 2989 19242 3155
rect -8216 -9304 -7656 -8744
<< metal3 >>
rect -15808 13017 20146 13500
rect -15808 12395 -4951 13017
rect -4393 13015 20146 13017
rect -4393 12395 16297 13015
rect -15808 12393 16297 12395
rect 16855 12393 20146 13015
rect -15808 12390 20146 12393
rect -4160 12388 20146 12390
rect 19496 4627 19672 12388
rect 15867 4609 16006 4614
rect 15867 4480 15872 4609
rect 16001 4480 16006 4609
rect 15867 4475 16006 4480
rect 18362 4609 18505 4614
rect 18362 4480 18367 4609
rect 18500 4480 18505 4609
rect 18362 4475 18505 4480
rect 15872 4096 16001 4475
rect 5539 3936 9821 3997
rect 15872 3968 16000 4096
rect 18369 4032 18498 4475
rect 19496 4461 19501 4627
rect 19620 4461 19672 4627
rect 19496 4456 19672 4461
rect 9979 3936 10437 3941
rect 5539 3488 9984 3936
rect 10432 3488 10437 3936
rect 5539 3427 9821 3488
rect 9979 3483 10437 3488
rect -8221 -8744 -7651 -8739
rect -8221 -9304 -8216 -8744
rect -7656 -9304 -7651 -8744
rect -8221 -12771 -7651 -9304
rect 5539 -12771 6109 3427
rect 15357 3145 15492 3459
rect 17854 3145 17989 3459
rect 19112 3155 19288 3160
rect 15351 3140 15497 3145
rect 15351 3005 15356 3140
rect 15492 3005 15497 3140
rect 15351 3000 15497 3005
rect 17848 3140 17994 3145
rect 17848 3005 17853 3140
rect 17989 3005 17994 3140
rect 17848 3000 17994 3005
rect 19112 2989 19117 3155
rect 19242 2989 19288 3155
rect 19112 -12771 19288 2989
rect -15837 -14109 20146 -12771
use JNW_VIS_ITIME  JNW_VIS_ITIME_0 ../JNW_GR02_SKY130A
timestamp 1744542523
transform 1 0 9649 0 1 12525
box -4353 -24590 9703 -1992
use JNW_VIS_TI  JNW_VIS_TI_0 ../JNW_GR02_SKY130A
timestamp 1744543763
transform 1 0 -5504 0 1 13448
box -9344 -19400 9900 -2398
use JNWTR_DFTSPCX1_CV  JNWTR_DFTSPCX1_CV_0 ../JNW_TR_SKY130A
timestamp 1744567443
transform 1 0 14690 0 1 3314
box -150 -120 2130 1080
use JNWTR_DFTSPCX1_CV  JNWTR_DFTSPCX1_CV_1
timestamp 1744567443
transform 1 0 17174 0 1 3320
box -150 -120 2130 1080
use JNW_VIS_TI  x2
timestamp 1744543763
transform 1 0 -5504 0 1 13448
box -9344 -19400 9900 -2398
use JNWTR_DFTSPCX1_CV  x3
timestamp 1744567443
transform 1 0 14690 0 1 3314
box -150 -120 2130 1080
use JNWTR_DFTSPCX1_CV  x4
timestamp 1744567443
transform 1 0 17174 0 1 3320
box -150 -120 2130 1080
<< labels >>
flabel metal3 -15836 12390 -4951 12958 0 FreeSans 1600 0 0 0 VDD_1V8
port 0 nsew
flabel metal3 -15168 448 -15040 576 0 FreeSans 1600 0 0 0 PWR_UP_1V8
port 11 nsew
flabel metal3 -15808 -13312 -15104 -13120 0 FreeSans 1600 0 0 0 VSS
port 1 nsew
flabel metal3 -15740 -10812 -13892 -10692 0 FreeSans 1600 0 0 0 CLK
port 21 nsew
flabel space 19968 4864 20096 4992 0 FreeSans 1600 0 0 0 VREF_OUT
port 22 nsew
<< properties >>
string FIXED_BBOX 0 0 22267 11539
<< end >>
