magic
tech sky130A
magscale 1 2
timestamp 1745877762
<< error_s >>
rect 17138 -15090 17148 -14990
rect 17218 -15090 17228 -14990
<< dnwell >>
rect 27560 -11240 34040 440
<< nwell >>
rect 27400 0 34400 1800
rect 27400 -10800 28000 0
rect 33600 -10800 34400 0
rect 27400 -11600 34400 -10800
<< nsubdiff >>
rect 30200 1200 31000 1400
rect 30200 1000 30400 1200
rect 30800 1000 31000 1200
rect 30200 800 31000 1000
<< nsubdiffcont >>
rect 30400 1000 30800 1200
<< locali >>
rect 30200 1200 31000 1400
rect 30200 1000 30400 1200
rect 30800 1000 31000 1200
rect 30200 800 31000 1000
rect 23804 -1010 37352 -1004
rect 23804 -1190 25078 -1010
rect 25258 -1190 37352 -1010
rect 23804 -1196 37352 -1190
rect 24688 -2224 24880 -1196
rect 26352 -2224 26544 -1196
rect 36456 -1458 36632 -1196
rect 29956 -1550 31306 -1490
rect 24688 -7250 24880 -4920
rect 26352 -5304 26544 -4872
rect 26096 -5496 26556 -5304
rect 26096 -5672 26288 -5496
rect 24688 -7430 24690 -7250
rect 24870 -7430 24880 -7250
rect 24688 -8644 24880 -7430
rect 26096 -8644 26288 -6884
rect 22220 -8836 26288 -8644
rect 24688 -10024 24880 -8836
rect 28976 -9260 29196 -1970
rect 29956 -2610 30016 -1550
rect 29416 -3130 29476 -2790
rect 30676 -3130 30736 -2810
rect 29416 -3142 30736 -3130
rect 29416 -3190 30676 -3142
rect 29956 -3970 30016 -3190
rect 29416 -4530 29476 -4230
rect 30676 -4530 30736 -4230
rect 29416 -4542 30736 -4530
rect 29416 -4590 30676 -4542
rect 29956 -5450 30016 -4590
rect 29416 -5970 29476 -5610
rect 30676 -5970 30736 -5630
rect 29416 -5982 30736 -5970
rect 29416 -6030 30676 -5982
rect 29956 -6870 30016 -6030
rect 29416 -7370 29476 -7030
rect 30676 -7370 30736 -7030
rect 29416 -7382 30736 -7370
rect 29416 -7430 30676 -7382
rect 29956 -8270 30016 -7430
rect 29416 -8770 29476 -8410
rect 30676 -8770 30736 -8410
rect 30976 -8720 31156 -1838
rect 31246 -5430 31306 -1550
rect 36456 -1622 36462 -1458
rect 36626 -1622 36632 -1458
rect 36456 -1628 36632 -1622
rect 36006 -2010 36216 -1950
rect 35180 -4898 35372 -2164
rect 36156 -2630 36216 -2010
rect 35616 -3250 35676 -2830
rect 36876 -3250 36936 -2810
rect 35616 -3310 36936 -3250
rect 36156 -3970 36216 -3310
rect 35616 -4490 35676 -4150
rect 36876 -4490 36936 -4170
rect 37160 -4436 37352 -1196
rect 35616 -4496 36936 -4490
rect 35616 -4544 36292 -4496
rect 36340 -4544 36936 -4496
rect 35616 -4550 36936 -4544
rect 35180 -5062 35194 -4898
rect 35358 -5062 35372 -4898
rect 31246 -5490 31998 -5430
rect 31246 -8770 31306 -5490
rect 29416 -8782 31306 -8770
rect 29416 -8830 30676 -8782
rect 30736 -8830 31306 -8782
rect 28976 -9390 29196 -9380
rect 35180 -10024 35372 -5062
rect 24688 -10216 35372 -10024
<< viali >>
rect 25078 -1190 25258 -1010
rect 24690 -7430 24870 -7250
rect 30976 -1838 31156 -1670
rect 30676 -3190 30736 -3142
rect 30676 -4590 30736 -4542
rect 30676 -6030 30736 -5982
rect 30676 -7430 30736 -7382
rect 36462 -1622 36626 -1458
rect 36292 -4544 36340 -4496
rect 35194 -5062 35358 -4898
rect 31998 -5490 32046 -5430
rect 30676 -8830 30736 -8782
rect 28976 -9380 29196 -9260
<< metal1 >>
rect 25072 -1010 25264 -998
rect 25072 -1190 25078 -1010
rect 25258 -1190 25264 -1010
rect 25072 -2356 25264 -1190
rect 36456 -1458 36632 -1446
rect 36456 -1622 36462 -1458
rect 36626 -1622 36632 -1458
rect 25968 -1670 31172 -1664
rect 25968 -1672 30976 -1670
rect 25968 -1848 30256 -1672
rect 30432 -1838 30976 -1672
rect 31156 -1838 31172 -1670
rect 36456 -1692 36632 -1622
rect 30432 -1848 31172 -1838
rect 25968 -1856 31172 -1848
rect 25968 -2316 26160 -1856
rect 36450 -1868 36456 -1692
rect 36632 -1868 36638 -1692
rect 24944 -3092 25008 -2708
rect 25072 -3176 25264 -2408
rect 30664 -3142 30748 -3136
rect 30664 -3190 30676 -3142
rect 30736 -3190 30748 -3142
rect 30664 -3196 30748 -3190
rect 30676 -3230 30736 -3196
rect 30676 -3296 30736 -3290
rect 24944 -3768 25008 -3468
rect 25968 -3640 26160 -3424
rect 25968 -3768 26496 -3640
rect 24944 -3832 26496 -3768
rect 24364 -4236 26156 -4044
rect 24364 -4312 24556 -4236
rect 23624 -4504 24556 -4312
rect 24944 -4412 25008 -4236
rect 25964 -4496 26156 -4236
rect 7904 -7156 8096 -5644
rect 24944 -6412 25008 -4968
rect 25072 -7244 25264 -4608
rect 26304 -5304 26496 -3832
rect 36286 -4496 36346 -4484
rect 30664 -4542 30748 -4536
rect 30664 -4590 30676 -4542
rect 30736 -4590 30748 -4542
rect 30664 -4596 30748 -4590
rect 36286 -4544 36292 -4496
rect 36340 -4544 36346 -4496
rect 30676 -4630 30736 -4596
rect 30676 -4696 30736 -4690
rect 35688 -4892 35864 -4886
rect 35182 -4898 35688 -4892
rect 35182 -5062 35194 -4898
rect 35358 -5062 35688 -4898
rect 35182 -5068 35688 -5062
rect 35688 -5074 35864 -5068
rect 25712 -5496 26496 -5304
rect 31992 -5430 32052 -5418
rect 36286 -5430 36346 -4544
rect 31992 -5490 31998 -5430
rect 32046 -5490 36346 -5430
rect 25712 -5704 25904 -5496
rect 31992 -5502 32052 -5490
rect 30664 -5982 30748 -5976
rect 30664 -6030 30676 -5982
rect 30736 -6030 30748 -5982
rect 30664 -6036 30748 -6030
rect 30676 -6070 30736 -6036
rect 30676 -6136 30736 -6130
rect 24678 -7250 25264 -7244
rect 24678 -7430 24690 -7250
rect 24870 -7430 25264 -7250
rect 24678 -7436 25264 -7430
rect 22888 -8092 23012 -8028
rect 22888 -8412 22952 -8092
rect 25712 -9245 25904 -6444
rect 30664 -7382 30748 -7376
rect 30664 -7430 30676 -7382
rect 30736 -7430 30748 -7382
rect 30664 -7436 30748 -7430
rect 30676 -7470 30736 -7436
rect 30676 -7536 30736 -7530
rect 30664 -8782 30748 -8776
rect 30664 -8830 30676 -8782
rect 30736 -8830 30748 -8782
rect 30664 -8836 30748 -8830
rect 30676 -8870 30736 -8836
rect 30676 -8936 30736 -8930
rect 25712 -9260 29421 -9245
rect 25712 -9376 28976 -9260
rect 25725 -9380 28976 -9376
rect 29196 -9380 29421 -9260
rect 25725 -9395 29421 -9380
rect 29571 -9395 29577 -9245
rect 20892 -15784 21084 -14744
rect 20684 -15976 21084 -15784
<< via1 >>
rect 30256 -1848 30432 -1672
rect 36456 -1868 36632 -1692
rect 30676 -3290 30736 -3230
rect 30676 -4690 30736 -4630
rect 35688 -5068 35864 -4892
rect 30676 -6130 30736 -6070
rect 30676 -7530 30736 -7470
rect 30676 -8930 30736 -8870
rect 29421 -9395 29571 -9245
<< metal2 >>
rect 30256 -1672 30432 -1666
rect 30256 -1957 30432 -1848
rect 36456 -1692 36632 -1686
rect 36456 -1937 36632 -1868
rect 30252 -2123 30261 -1957
rect 30427 -2123 30436 -1957
rect 36452 -2103 36461 -1937
rect 36627 -2103 36636 -1937
rect 36456 -2108 36632 -2103
rect 30256 -2128 30432 -2123
rect 30670 -3290 30676 -3230
rect 30736 -3290 30742 -3230
rect 30676 -3330 30736 -3290
rect 30517 -3390 30526 -3330
rect 30582 -3390 30736 -3330
rect 30670 -4690 30676 -4630
rect 30736 -4690 30742 -4630
rect 30676 -4730 30736 -4690
rect 30517 -4790 30526 -4730
rect 30582 -4790 30736 -4730
rect 35921 -4892 36087 -4888
rect 35682 -5068 35688 -4892
rect 35864 -4897 36092 -4892
rect 35864 -5063 35921 -4897
rect 36087 -5063 36092 -4897
rect 35864 -5068 36092 -5063
rect 35921 -5072 36087 -5068
rect 30670 -6130 30676 -6070
rect 30736 -6130 30742 -6070
rect 30676 -6170 30736 -6130
rect 30517 -6230 30526 -6170
rect 30582 -6230 30736 -6170
rect 30670 -7530 30676 -7470
rect 30736 -7530 30742 -7470
rect 30676 -7570 30736 -7530
rect 30517 -7630 30526 -7570
rect 30582 -7630 30736 -7570
rect 30670 -8930 30676 -8870
rect 30736 -8930 30742 -8870
rect 30676 -8970 30736 -8930
rect 30517 -9030 30526 -8970
rect 30582 -9030 30736 -8970
rect 29421 -9245 29571 -9239
rect 29571 -9395 29751 -9245
rect 29891 -9395 29900 -9245
rect 29421 -9401 29571 -9395
<< via2 >>
rect 30261 -2123 30427 -1957
rect 36461 -2103 36627 -1937
rect 30526 -3390 30582 -3330
rect 30526 -4790 30582 -4730
rect 35921 -5063 36087 -4897
rect 30526 -6230 30582 -6170
rect 30526 -7630 30582 -7570
rect 30526 -9030 30582 -8970
rect 29751 -9395 29891 -9245
<< metal3 >>
rect 36456 -1937 36632 -1932
rect 30256 -1957 30432 -1952
rect 30256 -2123 30261 -1957
rect 30427 -2123 30432 -1957
rect 29716 -9240 29892 -2692
rect 30256 -8652 30432 -2123
rect 36456 -2103 36461 -1937
rect 36627 -2103 36632 -1937
rect 30521 -3330 30587 -3325
rect 30521 -3390 30526 -3330
rect 30582 -3390 31886 -3330
rect 30521 -3395 30587 -3390
rect 30521 -4730 30587 -4725
rect 30521 -4790 30526 -4730
rect 30582 -4790 31906 -4730
rect 30521 -4795 30587 -4790
rect 35916 -4897 36092 -2852
rect 36456 -3888 36632 -2103
rect 35916 -5063 35921 -4897
rect 36087 -5063 36092 -4897
rect 35916 -5068 36092 -5063
rect 30521 -6170 30587 -6165
rect 30521 -6230 30526 -6170
rect 30582 -6230 32006 -6170
rect 30521 -6235 30587 -6230
rect 30521 -7570 30587 -7565
rect 30521 -7630 30526 -7570
rect 30582 -7630 31966 -7570
rect 30521 -7635 30587 -7630
rect 30521 -8970 30587 -8965
rect 30521 -9030 30526 -8970
rect 30582 -9030 32026 -8970
rect 30521 -9035 30587 -9030
rect 29716 -9245 29896 -9240
rect 29716 -9395 29751 -9245
rect 29891 -9395 29983 -9245
rect 30131 -9395 30137 -9245
rect 29716 -9400 29896 -9395
rect 29716 -9408 29892 -9400
<< via3 >>
rect 29983 -9395 30131 -9245
<< metal4 >>
rect 29982 -9245 30132 -9244
rect 32321 -9245 32471 -3695
rect 29982 -9395 29983 -9245
rect 30131 -9395 32471 -9245
rect 29982 -9396 30132 -9395
rect 17030 -15090 17330 -14990
use JNWTR_CAPX1  JNWTR_CAPX1_0 ../JNW_TR_SKY130A
timestamp 1745877762
transform 0 1 31636 1 0 -9720
box 0 0 1080 1080
use JNWTR_IVX4_CV  JNWTR_IVX4_CV_0 ../JNW_TR_SKY130A
timestamp 1745877762
transform 1 0 29086 0 1 -8680
box -150 -120 2130 920
use JNWTR_IVX4_CV  JNWTR_IVX4_CV_1
timestamp 1745877762
transform 1 0 29086 0 1 -4380
box -150 -120 2130 920
use JNWTR_IVX4_CV  JNWTR_IVX4_CV_2
timestamp 1745877762
transform 1 0 29086 0 1 -7180
box -150 -120 2130 920
use JNWTR_IVX4_CV  JNWTR_IVX4_CV_3
timestamp 1745877762
transform 1 0 29086 0 1 -5880
box -150 -120 2130 920
use JNWTR_IVX4_CV  JNWTR_IVX4_CV_4
timestamp 1745877762
transform 1 0 29086 0 1 -2980
box -150 -120 2130 920
use JNW_VIS_TI  x2 ../JNW_GR02_SKY130A
timestamp 1745877762
transform 1 0 14388 0 1 1400
box -9344 -19400 9900 -2398
use JNWTR_CAPX1  x7
timestamp 1745877762
transform 0 -1 32716 1 0 -3800
box 0 0 1080 1080
use JNWATR_NCH_8C1F2  x8 ../JNW_ATR_SKY130A
timestamp 1745877762
transform 1 0 24784 0 1 -7072
box -184 -128 1592 928
use JNWATR_NCH_12C1F2  x9 ../JNW_ATR_SKY130A
timestamp 1745877762
transform 1 0 24784 0 1 -5072
box -184 -128 1848 928
use JNWTR_IVX4_CV  x10
timestamp 1745877762
transform 1 0 35286 0 1 -3080
box -150 -120 2130 920
use JNWATR_NCH_8C1F2  x11
timestamp 1745877762
transform 1 0 24784 0 1 -6272
box -184 -128 1592 928
use JNWATR_PCH_12C1F2  x12 ../JNW_ATR_SKY130A
timestamp 1745877762
transform 1 0 24784 0 1 -3672
box -184 -128 1848 928
use JNWATR_PCH_12C1F2  x13
timestamp 1745877762
transform 1 0 24784 0 1 -2872
box -184 -128 1848 928
use JNWTR_IVX4_CV  x14
timestamp 1745877762
transform 1 0 35286 0 1 -4420
box -150 -120 2130 920
use JNWTR_CAPX1  x15
timestamp 1745877762
transform 0 -1 32716 1 0 -5300
box 0 0 1080 1080
use JNWTR_CAPX1  x16
timestamp 1745877762
transform 0 -1 32716 1 0 -6800
box 0 0 1080 1080
use JNWTR_CAPX1  x17
timestamp 1745877762
transform 0 -1 32716 1 0 -8300
box 0 0 1080 1080
<< labels >>
flabel locali 24688 -10216 26686 -10024 0 FreeSans 1600 0 0 0 VSS
port 0 nsew
flabel metal1 22948 -8092 23012 -8028 0 FreeSans 1600 0 0 0 PWR_UP
port 2 nsew
flabel locali 36006 -2010 36066 -1950 0 FreeSans 1600 0 0 0 VOUT
port 1 nsew
flabel metal1 7904 -5836 8096 -5644 0 FreeSans 1600 0 0 0 VREF
port 4 nsew
flabel locali 29460 -1196 29652 -1004 0 FreeSans 1600 0 0 0 VDD
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 34124 12080
<< end >>
